* Design:	NAND2x1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2x1_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00570454f
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00471464f
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%A VSS 19 3 4 5 1
c1 1 VSS 0.00708684f
c2 3 VSS 0.0431806f
c3 4 VSS 0.080425f
c4 5 VSS 0.00806292f
c5 6 VSS 0.0135161f
c6 7 VSS 0.00361733f
c7 8 VSS 0.00249676f
r1 6 8 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1350
r2 5 8 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1160 $X2=0.0270 $Y2=0.1350
r3 8 21 1.38478 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0380 $Y2=0.1350
r4 4 17 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1345
r5 19 7 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0505 $Y2=0.1350
r6 7 21 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0505
+ $Y=0.1350 $X2=0.0380 $Y2=0.1350
r7 15 17 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1345 $X2=0.1350 $Y2=0.1345
r8 14 15 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1345 $X2=0.1225 $Y2=0.1345
r9 13 14 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1345 $X2=0.1080 $Y2=0.1345
r10 1 9 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1345 $X2=0.0850 $Y2=0.1345
r11 1 10 2.09261 $w=2.04231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0750 $Y=0.1345 $X2=0.0685 $Y2=0.1345
r12 19 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1345
r13 3 9 1.73446 $w=1.505e-07 $l=4.03113e-09 $layer=LIG $thickness=5.3e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0850 $Y2=0.1345
r14 3 10 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1345
r15 3 13 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1345
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00543988f
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00463639f
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%B VSS 18 3 4 1 5
c1 1 VSS 0.0112506f
c2 3 VSS 0.0472567f
c3 4 VSS 0.00984508f
c4 5 VSS 0.0057051f
r1 18 17 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1520 $X2=0.2430 $Y2=0.1477
r2 5 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r3 5 17 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1477
r4 4 13 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 10 12 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2335 $Y2=0.1350
r7 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2305 $Y2=0.1350
r8 8 9 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2015
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r9 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r10 1 7 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r11 1 8 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r12 3 7 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r13 3 8 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%NET16 VSS 15 27 28 30 1 2 13 10 11 3 12
c1 1 VSS 0.0080921f
c2 2 VSS 0.00752539f
c3 3 VSS 0.00533166f
c4 10 VSS 0.00342352f
c5 11 VSS 0.00337042f
c6 12 VSS 0.00223029f
c7 13 VSS 0.0220178f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r2 30 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r3 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r4 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r6 27 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r7 3 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r8 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r9 22 23 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r10 21 22 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1865
+ $Y=0.0360 $X2=0.2315 $Y2=0.0360
r11 20 21 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1865 $Y2=0.0360
r12 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r13 18 19 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0890
+ $Y=0.0360 $X2=0.1235 $Y2=0.0360
r14 17 18 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0735
+ $Y=0.0360 $X2=0.0890 $Y2=0.0360
r15 16 17 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0735 $Y2=0.0360
r16 13 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r17 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r18 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r19 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r20 1 10 1e-05
.ends

.subckt PM_NAND2x1_ASAP7_75t_R%Y VSS 29 19 22 40 42 13 1 11 12 14 2 3 15 10
c1 1 VSS 0.00841902f
c2 2 VSS 0.00294319f
c3 3 VSS 0.00787406f
c4 10 VSS 0.00211307f
c5 11 VSS 0.00354207f
c6 12 VSS 0.00345751f
c7 13 VSS 0.0191991f
c8 14 VSS 0.00082208f
c9 15 VSS 0.00233706f
c10 16 VSS 0.000770033f
c11 17 VSS 0.00298135f
r1 42 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 11 41 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r4 40 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 1 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r7 37 38 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1595 $Y2=0.2340
r8 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r9 33 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r10 33 38 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.1595 $Y2=0.2340
r11 32 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r12 13 17 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2970 $Y2=0.2340
r13 13 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r14 17 31 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2970 $Y2=0.2125
r15 30 31 9.26929 $w=1.3e-08 $l=3.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1727 $X2=0.2970 $Y2=0.2125
r16 29 30 6.47102 $w=1.3e-08 $l=2.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1450 $X2=0.2970 $Y2=0.1727
r17 29 28 4.6055 $w=1.3e-08 $l=1.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1450 $X2=0.2970 $Y2=0.1252
r18 15 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0935 $X2=0.2970 $Y2=0.0720
r19 15 28 7.40377 $w=1.3e-08 $l=3.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0935 $X2=0.2970 $Y2=0.1252
r20 16 27 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0720 $X2=0.2860 $Y2=0.0720
r21 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.0720 $X2=0.2860 $Y2=0.0720
r22 25 26 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0720 $X2=0.2680 $Y2=0.0720
r23 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r24 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.2295 $Y2=0.0720
r25 14 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r26 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r27 22 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r28 20 21 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r29 2 20 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0675 $X2=0.2260 $Y2=0.0675
r30 10 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r31 19 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r32 1 11 1e-05
.ends


*
.SUBCKT NAND2x1_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM3@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NAND2x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2x1_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2x1_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM3_g 0.00243823f
cc_2 N_noxref_7_1 N_NET16_10 0.0363555f
x_PM_NAND2x1_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2x1_ASAP7_75t_R%noxref_8
cc_3 N_noxref_8_1 N_MM3_g 0.0104487f
cc_4 N_noxref_8_1 N_NET16_10 0.000601385f
cc_5 N_noxref_8_1 N_Y_11 0.000624583f
cc_6 N_noxref_8_1 N_noxref_7_1 0.00191604f
x_PM_NAND2x1_ASAP7_75t_R%A VSS A N_MM3_g N_MM3@2_g N_A_5 N_A_1
+ PM_NAND2x1_ASAP7_75t_R%A
x_PM_NAND2x1_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2x1_ASAP7_75t_R%noxref_9
cc_7 N_noxref_9_1 N_MM2@2_g 0.00166953f
cc_8 N_noxref_9_1 N_NET16_12 0.0364845f
cc_9 N_noxref_9_1 N_Y_10 0.000787723f
x_PM_NAND2x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2x1_ASAP7_75t_R%noxref_10
cc_10 N_noxref_10_1 N_MM2@2_g 0.00919382f
cc_11 N_noxref_10_1 N_NET16_12 0.000643758f
cc_12 N_noxref_10_1 N_Y_12 0.00185021f
cc_13 N_noxref_10_1 N_noxref_9_1 0.00193489f
x_PM_NAND2x1_ASAP7_75t_R%B VSS B N_MM2_g N_MM2@2_g N_B_1 N_B_5
+ PM_NAND2x1_ASAP7_75t_R%B
cc_14 N_MM2_g N_MM3@2_g 0.00476266f
x_PM_NAND2x1_ASAP7_75t_R%NET16 VSS N_MM3_d N_MM3@2_d N_MM2_s N_MM2@2_s
+ N_NET16_1 N_NET16_2 N_NET16_13 N_NET16_10 N_NET16_11 N_NET16_3 N_NET16_12
+ PM_NAND2x1_ASAP7_75t_R%NET16
cc_15 N_NET16_1 N_MM3_g 0.00269925f
cc_16 N_NET16_2 N_MM3@2_g 0.000884991f
cc_17 N_NET16_13 N_MM3@2_g 0.00131002f
cc_18 N_NET16_13 N_A_5 0.00169345f
cc_19 N_NET16_10 N_A_1 0.00214173f
cc_20 N_NET16_11 N_MM3@2_g 0.0333808f
cc_21 N_NET16_10 N_MM3_g 0.0357728f
cc_22 N_NET16_2 N_MM2@2_g 0.000877321f
cc_23 N_NET16_3 N_MM2@2_g 0.00109033f
cc_24 N_NET16_12 N_B_1 0.00169018f
cc_25 N_NET16_11 N_MM2_g 0.0335036f
cc_26 N_NET16_12 N_MM2@2_g 0.0358182f
x_PM_NAND2x1_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM2@2_d N_MM1_d N_MM0_d N_Y_13 N_Y_1
+ N_Y_11 N_Y_12 N_Y_14 N_Y_2 N_Y_3 N_Y_15 N_Y_10 PM_NAND2x1_ASAP7_75t_R%Y
cc_27 N_Y_13 N_MM3@2_g 0.000764315f
cc_28 N_Y_1 N_MM3@2_g 0.00263063f
cc_29 N_Y_11 N_A_1 0.00266984f
cc_30 N_Y_11 N_MM3_g 0.0191786f
cc_31 N_Y_11 N_MM3@2_g 0.0542245f
cc_32 N_Y_12 N_MM2_g 0.012028f
cc_33 N_Y_14 N_B_5 0.0012637f
cc_34 N_Y_13 N_B_5 0.00147115f
cc_35 N_Y_2 N_MM2@2_g 0.00189817f
cc_36 N_Y_3 N_MM2@2_g 0.00268656f
cc_37 N_Y_12 N_B_1 0.00477819f
cc_38 N_Y_15 N_B_5 0.00765093f
cc_39 N_Y_12 N_MM2@2_g 0.0212458f
cc_40 N_Y_10 N_MM2_g 0.0374567f
cc_41 N_Y_10 N_MM2@2_g 0.0707371f
cc_42 N_Y_14 N_NET16_3 0.000667538f
cc_43 N_Y_10 N_NET16_12 0.0018262f
cc_44 N_Y_15 N_NET16_3 0.000735448f
cc_45 N_Y_2 N_NET16_13 0.000818119f
cc_46 N_Y_2 N_NET16_2 0.00151578f
cc_47 N_Y_2 N_NET16_3 0.005261f
cc_48 N_Y_14 N_NET16_13 0.0102134f
*END of NAND2x1_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND2x1p5_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2x1p5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2x1p5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2x1p5_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0420017f
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00519099f
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00534879f
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00467014f
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%A VSS 26 3 4 5 1 8
c1 1 VSS 0.0129976f
c2 3 VSS 0.043484f
c3 4 VSS 0.0799217f
c4 5 VSS 0.0803353f
c5 6 VSS 0.0177448f
c6 7 VSS 0.0170548f
c7 8 VSS 0.00375127f
c8 9 VSS 0.00326603f
r1 7 9 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1350
r2 6 9 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.1350
r3 5 24 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1345
r4 4 18 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1345
r5 26 8 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0485 $Y2=0.1350
r6 8 9 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0485
+ $Y=0.1350 $X2=0.0270 $Y2=0.1350
r7 22 24 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1345 $X2=0.1890 $Y2=0.1345
r8 21 22 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1345 $X2=0.1765 $Y2=0.1345
r9 19 21 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1345 $X2=0.1620 $Y2=0.1345
r10 18 19 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1345 $X2=0.1475 $Y2=0.1345
r11 16 18 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1345 $X2=0.1350 $Y2=0.1345
r12 15 16 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1345 $X2=0.1225 $Y2=0.1345
r13 14 15 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1345 $X2=0.1080 $Y2=0.1345
r14 1 10 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1345 $X2=0.0850 $Y2=0.1345
r15 1 11 2.09261 $w=2.04231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0750 $Y=0.1345 $X2=0.0685 $Y2=0.1345
r16 26 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1345
r17 3 10 1.73446 $w=1.505e-07 $l=4.03113e-09 $layer=LIG $thickness=5.3e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0850 $Y2=0.1345
r18 3 11 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1345
r19 3 14 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1345
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%NET16 VSS 17 20 35 36 38 41 1 11 12 13 14 3 15
+ 2
c1 1 VSS 0.00999435f
c2 2 VSS 0.00749886f
c3 3 VSS 0.00285341f
c4 11 VSS 0.00440823f
c5 12 VSS 0.00319671f
c6 13 VSS 0.00208068f
c7 14 VSS 0.0121628f
c8 15 VSS 0.00163327f
r1 41 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r2 39 40 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r3 3 39 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0675 $X2=0.3340 $Y2=0.0675
r4 13 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 38 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0720
r7 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r8 2 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r9 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r10 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r11 30 31 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2880
+ $Y=0.0720 $X2=0.3240 $Y2=0.0720
r12 29 30 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2590
+ $Y=0.0720 $X2=0.2880 $Y2=0.0720
r13 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2410
+ $Y=0.0720 $X2=0.2590 $Y2=0.0720
r14 27 28 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.2410 $Y2=0.0720
r15 15 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r16 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r17 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r18 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r19 24 25 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1730
+ $Y=0.0360 $X2=0.2045 $Y2=0.0360
r20 23 24 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1730 $Y2=0.0360
r21 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r22 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r23 14 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r24 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r25 20 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r26 1 19 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r27 16 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.0675 $X2=0.1100 $Y2=0.0675
r28 11 16 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.0980 $Y2=0.0675
r29 17 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%B VSS 30 3 4 5 7 9 8 6 1
c1 1 VSS 0.0139496f
c2 3 VSS 0.0467974f
c3 4 VSS 0.0463455f
c4 5 VSS 0.00940555f
c5 6 VSS 0.00576779f
c6 7 VSS 0.00578127f
c7 8 VSS 0.00631165f
c8 9 VSS 0.00432627f
r1 7 31 6.91198 $w=1.35906e-08 $l=3.18e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1720 $X2=0.1350 $Y2=0.1402
r2 6 9 5.73148 $w=1.38716e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1307
r3 30 31 0.433689 $w=1.8e-08 $l=4.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.1402
r4 30 9 0.535733 $w=1.8e-08 $l=5.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.1307
r5 5 24 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 4 18 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r7 30 28 6.81353 $w=1.01579e-08 $l=3.80132e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1360 $X2=0.1730 $Y2=0.1350
r8 8 26 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r9 8 28 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1350 $X2=0.1730 $Y2=0.1350
r10 22 24 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r11 21 22 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r12 19 21 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r13 18 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r14 16 18 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r15 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r17 12 14 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2525 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r18 11 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2525 $Y2=0.1350
r19 11 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r20 1 11 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r21 1 13 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2325 $Y2=0.1350
r22 3 11 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r23 3 13 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r24 3 14 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NAND2x1p5_ASAP7_75t_R%Y VSS 39 27 30 43 55 58 59 61 2 21 1 18 19 3
+ 17 23 5 20 4 16 22
c1 1 VSS 0.00795189f
c2 2 VSS 0.00908914f
c3 3 VSS 0.00452356f
c4 4 VSS 0.00780471f
c5 5 VSS 0.00513475f
c6 16 VSS 0.00218936f
c7 17 VSS 0.00232217f
c8 18 VSS 0.00349782f
c9 19 VSS 0.00415321f
c10 20 VSS 0.0034756f
c11 21 VSS 0.0294951f
c12 22 VSS 0.0113003f
c13 23 VSS 0.00346042f
c14 24 VSS 0.00283669f
c15 25 VSS 0.00297196f
r1 61 60 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 18 60 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r4 2 57 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r5 19 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r6 58 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r7 20 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r8 55 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r9 1 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r10 2 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r11 4 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r12 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r13 50 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r14 48 49 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2410 $Y2=0.2340
r15 47 48 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r16 47 50 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 45 46 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3355 $Y2=0.2340
r18 44 45 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r19 44 49 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.2340 $X2=0.2410 $Y2=0.2340
r20 21 25 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3670 $Y=0.2340 $X2=0.4050 $Y2=0.2340
r21 21 46 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.2340 $X2=0.3355 $Y2=0.2340
r22 25 41 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.4050 $Y2=0.2125
r23 17 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3760 $Y2=0.0675
r24 43 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r25 40 41 9.26929 $w=1.3e-08 $l=3.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1727 $X2=0.4050 $Y2=0.2125
r26 39 40 6.47102 $w=1.3e-08 $l=2.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1450 $X2=0.4050 $Y2=0.1727
r27 39 38 0.174892 $w=1.3e-08 $l=8e-10 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1450 $X2=0.4050 $Y2=0.1442
r28 37 38 2.15701 $w=1.3e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1442
r29 36 37 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1035 $X2=0.4050 $Y2=0.1350
r30 35 36 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0720 $X2=0.4050 $Y2=0.1035
r31 23 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0360
r32 23 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0720
r33 5 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r34 24 34 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3915 $Y2=0.0360
r35 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r36 32 33 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r37 31 32 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3535 $Y2=0.0360
r38 22 31 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3085 $Y2=0.0360
r39 3 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r40 30 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r41 3 29 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r42 26 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2600 $Y=0.0675 $X2=0.2720 $Y2=0.0675
r43 16 26 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2600 $Y2=0.0675
r44 27 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r45 1 18 1e-05
.ends


*
.SUBCKT NAND2x1p5_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@3 N_MM3@3_d N_MM3@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM3@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@3 N_MM2@3_d N_MM2@3_g N_MM2@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 N_MM1@2_d N_MM2@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NAND2x1p5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2x1p5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2x1p5_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2x1p5_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM3_g 0.00253354f
x_PM_NAND2x1p5_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2x1p5_ASAP7_75t_R%noxref_9
cc_2 N_noxref_9_1 N_MM2@2_g 0.00163091f
cc_3 N_noxref_9_1 N_Y_17 0.0376033f
x_PM_NAND2x1p5_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2x1p5_ASAP7_75t_R%noxref_8
cc_4 N_noxref_8_1 N_MM3_g 0.0105162f
cc_5 N_noxref_8_1 N_Y_18 0.000609858f
cc_6 N_noxref_8_1 N_noxref_7_1 0.00192564f
x_PM_NAND2x1p5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2x1p5_ASAP7_75t_R%noxref_10
cc_7 N_noxref_10_1 N_MM2@2_g 0.00902823f
cc_8 N_noxref_10_1 N_Y_20 0.00262698f
cc_9 N_noxref_10_1 N_noxref_9_1 0.00193469f
x_PM_NAND2x1p5_ASAP7_75t_R%A VSS A N_MM3_g N_MM3@3_g N_MM3@2_g N_A_1 N_A_8
+ PM_NAND2x1p5_ASAP7_75t_R%A
x_PM_NAND2x1p5_ASAP7_75t_R%NET16 VSS N_MM3_d N_MM3@3_d N_MM3@2_d N_MM2_s
+ N_MM2@3_s N_MM2@2_s N_NET16_1 N_NET16_11 N_NET16_12 N_NET16_13 N_NET16_14
+ N_NET16_3 N_NET16_15 N_NET16_2 PM_NAND2x1p5_ASAP7_75t_R%NET16
cc_10 N_NET16_1 N_MM3@3_g 0.00203759f
cc_11 N_NET16_11 N_A_1 0.00313426f
cc_12 N_NET16_12 N_MM3@2_g 0.0328978f
cc_13 N_NET16_11 N_MM3_g 0.0181182f
cc_14 N_NET16_11 N_MM3@3_g 0.0509859f
cc_15 N_NET16_13 N_MM2_g 0.00101922f
cc_16 N_NET16_14 N_B_6 0.00138364f
cc_17 N_NET16_3 N_MM2@2_g 0.00168274f
cc_18 N_NET16_1 N_B_6 0.00244367f
cc_19 N_NET16_13 N_B_1 0.0031724f
cc_20 N_NET16_15 N_B_8 0.00338954f
cc_21 N_NET16_12 N_MM2_g 0.0329442f
cc_22 N_NET16_13 N_MM2@3_g 0.0181163f
cc_23 N_NET16_13 N_MM2@2_g 0.0499429f
x_PM_NAND2x1p5_ASAP7_75t_R%B VSS B N_MM2_g N_MM2@3_g N_MM2@2_g N_B_7 N_B_9
+ N_B_8 N_B_6 N_B_1 PM_NAND2x1p5_ASAP7_75t_R%B
cc_24 N_B_7 N_A_1 0.000946066f
cc_25 N_B_9 N_A_8 0.000946315f
cc_26 N_B_8 N_A_1 0.000965262f
cc_27 N_B_9 N_A_1 0.00252523f
cc_28 N_MM2_g N_MM3@2_g 0.00784236f
x_PM_NAND2x1p5_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM2@3_d N_MM2@2_d N_MM1@2_d
+ N_MM0@2_d N_MM1_d N_MM0_d N_Y_2 N_Y_21 N_Y_1 N_Y_18 N_Y_19 N_Y_3 N_Y_17
+ N_Y_23 N_Y_5 N_Y_20 N_Y_4 N_Y_16 N_Y_22 PM_NAND2x1p5_ASAP7_75t_R%Y
cc_29 N_Y_2 N_MM3@3_g 0.000356419f
cc_30 N_Y_21 N_MM3@3_g 0.00121809f
cc_31 N_Y_1 N_MM3@3_g 0.00252008f
cc_32 N_Y_18 N_A_1 0.00253843f
cc_33 N_Y_19 N_MM3@2_g 0.0242546f
cc_34 N_Y_18 N_MM3_g 0.0191027f
cc_35 N_Y_18 N_MM3@3_g 0.0531528f
cc_36 N_Y_3 N_MM2@3_g 0.00234785f
cc_37 N_Y_17 N_MM2@3_g 0.000452218f
cc_38 N_Y_2 N_MM2@3_g 0.000610012f
cc_39 N_Y_23 N_B_1 0.000789928f
cc_40 N_Y_5 N_MM2@2_g 0.000889309f
cc_41 N_Y_20 N_MM2@3_g 0.0119472f
cc_42 N_Y_2 N_B_8 0.00126132f
cc_43 N_Y_4 N_MM2@2_g 0.00223624f
cc_44 N_Y_21 N_B_8 0.00237987f
cc_45 N_Y_1 N_B_7 0.00241466f
cc_46 N_Y_19 N_MM2_g 0.0108177f
cc_47 N_Y_20 N_B_1 0.00636473f
cc_48 N_Y_17 N_MM2@2_g 0.053476f
cc_49 N_Y_20 N_MM2@2_g 0.0211903f
cc_50 N_Y_16 N_MM2_g 0.0321868f
cc_51 N_Y_16 N_MM2@3_g 0.0692846f
cc_52 N_Y_3 N_NET16_15 0.00112045f
cc_53 N_Y_16 N_NET16_15 0.000557273f
cc_54 N_Y_17 N_NET16_15 0.00056165f
cc_55 N_Y_23 N_NET16_15 0.000652587f
cc_56 N_Y_22 N_NET16_3 0.000922673f
cc_57 N_Y_17 N_NET16_13 0.00111274f
cc_58 N_Y_16 N_NET16_13 0.00111627f
cc_59 N_Y_3 N_NET16_2 0.00117088f
cc_60 N_Y_3 N_NET16_3 0.00316752f
cc_61 N_Y_5 N_NET16_3 0.00432892f
cc_62 N_Y_22 N_NET16_15 0.0106018f
*END of NAND2x1p5_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND2x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2x2_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00589468f
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00584711f
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0046437f
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00462958f
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%A VSS 30 3 4 5 6 7 1 8
c1 1 VSS 0.02095f
c2 3 VSS 0.0843799f
c3 4 VSS 0.0472281f
c4 5 VSS 0.0472324f
c5 6 VSS 0.0843506f
c6 7 VSS 0.00519215f
c7 8 VSS 0.00474435f
r1 8 32 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2700 $Y2=0.1830
r2 3 26 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1345
r3 4 20 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1345
r4 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1605 $X2=0.2700 $Y2=0.1830
r5 30 31 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2700 $Y2=0.1605
r6 30 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2700 $Y2=0.1215
r7 7 29 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1115 $X2=0.2700 $Y2=0.1215
r8 5 14 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1345
r9 24 26 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1345 $X2=0.1890 $Y2=0.1345
r10 23 24 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1345 $X2=0.2015 $Y2=0.1345
r11 21 23 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1345 $X2=0.2160 $Y2=0.1345
r12 20 21 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1345 $X2=0.2305 $Y2=0.1345
r13 18 20 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1345 $X2=0.2430 $Y2=0.1345
r14 17 18 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1345 $X2=0.2555 $Y2=0.1345
r15 30 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2700 $Y=0.1350
+ $X2=0.2700 $Y2=0.1345
r16 15 17 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1345 $X2=0.2700 $Y2=0.1345
r17 14 15 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1345 $X2=0.2845 $Y2=0.1345
r18 12 14 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1345 $X2=0.2970 $Y2=0.1345
r19 11 12 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1345 $X2=0.3095 $Y2=0.1345
r20 10 11 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1345 $X2=0.3240 $Y2=0.1345
r21 6 1 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1345
r22 1 10 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1345 $X2=0.3385 $Y2=0.1345
r23 1 28 2.59554 $w=2.2681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1345 $X2=0.3615 $Y2=0.1345
r24 6 10 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3385 $Y2=0.1345
r25 6 28 0.54388 $w=2.16967e-07 $l=1.05119e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.3510 $Y=0.1350 $X2=0.3615 $Y2=0.1345
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%B VSS 34 5 6 7 8 12 1 2 10 19 14 21 16 13 11 18
+ 20 17 22 9 15
c1 1 VSS 0.00658975f
c2 2 VSS 0.00660571f
c3 5 VSS 0.00757088f
c4 6 VSS 0.0447943f
c5 7 VSS 0.0447975f
c6 8 VSS 0.00755902f
c7 9 VSS 0.00294244f
c8 10 VSS 0.00371401f
c9 11 VSS 0.00285012f
c10 12 VSS 0.00455022f
c11 13 VSS 0.00285497f
c12 14 VSS 0.00370543f
c13 15 VSS 0.00301235f
c14 16 VSS 0.00250433f
c15 17 VSS 0.0030803f
c16 18 VSS 0.00299739f
c17 19 VSS 0.00284424f
c18 20 VSS 0.00302621f
c19 21 VSS 0.00288828f
c20 22 VSS 0.00249638f
r1 7 55 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r2 8 48 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r3 53 55 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 52 53 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r5 50 52 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r6 2 48 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r7 2 50 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4465 $Y2=0.1350
r8 46 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r9 15 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1215 $X2=0.4590 $Y2=0.1350
r10 15 22 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1215 $X2=0.4590 $Y2=0.1080
r11 22 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1080 $X2=0.4340 $Y2=0.1080
r12 14 21 9.45156 $w=1.34118e-08 $l=4.83141e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3790 $Y=0.1080 $X2=0.3310 $Y2=0.1025
r13 14 45 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3790
+ $Y=0.1080 $X2=0.4340 $Y2=0.1080
r14 13 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.0900 $X2=0.3310 $Y2=0.0720
r15 13 21 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3310 $Y=0.0900 $X2=0.3310 $Y2=0.1025
r16 20 43 5.46317 $w=1.44754e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3310 $Y=0.0720 $X2=0.3005 $Y2=0.0720
r17 42 43 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0720 $X2=0.3005 $Y2=0.0720
r18 41 42 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2515
+ $Y=0.0720 $X2=0.2700 $Y2=0.0720
r19 12 18 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2300 $Y=0.0720 $X2=0.2090 $Y2=0.0720
r20 12 41 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2300
+ $Y=0.0720 $X2=0.2515 $Y2=0.0720
r21 11 19 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2090 $Y=0.0900 $X2=0.2090 $Y2=0.1025
r22 11 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.0900 $X2=0.2090 $Y2=0.0720
r23 19 39 9.45156 $w=1.34118e-08 $l=4.83141e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2090 $Y=0.1025 $X2=0.1610 $Y2=0.1080
r24 38 39 10.6101 $w=1.3e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1155
+ $Y=0.1080 $X2=0.1610 $Y2=0.1080
r25 10 16 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0995 $Y=0.1080 $X2=0.0810 $Y2=0.1080
r26 10 38 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0995
+ $Y=0.1080 $X2=0.1155 $Y2=0.1080
r27 17 35 5.17411 $w=1.46514e-08 $l=2.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1980 $X2=0.0810 $Y2=0.1707
r28 6 30 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r29 34 35 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1520 $X2=0.0810 $Y2=0.1707
r30 34 33 0.991057 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1520 $X2=0.0810 $Y2=0.1477
r31 32 33 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1477
r32 9 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1215 $X2=0.0810 $Y2=0.1350
r33 9 16 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1215 $X2=0.0810 $Y2=0.1080
r34 28 30 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r35 27 28 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r36 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r37 24 26 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r38 23 24 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r39 23 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r40 1 23 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r41 1 25 0.721303 $w=1.75333e-08 $l=1.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0715 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r42 5 23 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r43 5 25 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r44 5 26 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%NET16 VSS 23 40 41 44 45 48 49 51 16 21 1 5 3 17
+ 20 19 4 2 18
c1 1 VSS 0.00524237f
c2 2 VSS 0.00708705f
c3 3 VSS 0.00909804f
c4 4 VSS 0.00724924f
c5 5 VSS 0.0052577f
c6 16 VSS 0.00221228f
c7 17 VSS 0.00332719f
c8 18 VSS 0.00435975f
c9 19 VSS 0.0033339f
c10 20 VSS 0.00221068f
c11 21 VSS 0.0386435f
r1 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 51 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r4 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r5 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r6 48 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r7 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r8 3 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r9 18 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r10 44 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r11 41 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r12 2 39 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r13 17 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r14 40 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r15 5 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r16 4 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r17 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r18 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r19 35 36 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r20 34 35 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4025
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r21 33 34 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4025 $Y2=0.0360
r22 32 33 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3545
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r23 31 32 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3095
+ $Y=0.0360 $X2=0.3545 $Y2=0.0360
r24 30 31 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3095 $Y2=0.0360
r25 29 30 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2305
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r26 28 29 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1855
+ $Y=0.0360 $X2=0.2305 $Y2=0.0360
r27 27 28 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1855 $Y2=0.0360
r28 26 27 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1375
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r29 25 26 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0925
+ $Y=0.0360 $X2=0.1375 $Y2=0.0360
r30 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0925 $Y2=0.0360
r31 21 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r32 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r33 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r34 16 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r35 1 16 1e-05
.ends

.subckt PM_NAND2x2_ASAP7_75t_R%Y VSS 73 35 38 63 65 67 69 81 84 4 3 2 1 5 6 19
+ 24 21 26 28 27 25 29 20 23 22 32 30
c1 1 VSS 0.00289613f
c2 2 VSS 0.0076679f
c3 3 VSS 0.00755026f
c4 4 VSS 0.00770526f
c5 5 VSS 0.00290957f
c6 6 VSS 0.00770222f
c7 19 VSS 0.00211925f
c8 20 VSS 0.00211804f
c9 21 VSS 0.00346096f
c10 22 VSS 0.00347009f
c11 23 VSS 0.0034671f
c12 24 VSS 0.00345054f
c13 25 VSS 0.00227335f
c14 26 VSS 0.000645577f
c15 27 VSS 0.0392909f
c16 28 VSS 0.000697926f
c17 29 VSS 0.00236962f
c18 30 VSS 0.000792149f
c19 31 VSS 0.00283177f
c20 32 VSS 0.000792332f
c21 33 VSS 0.00298087f
r1 84 83 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r2 82 83 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r3 5 82 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0675 $X2=0.4420 $Y2=0.0675
r4 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r5 81 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r6 5 78 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0720
r7 78 79 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0720 $X2=0.4545 $Y2=0.0720
r8 76 79 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.0720 $X2=0.4545 $Y2=0.0720
r9 28 32 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5020 $Y=0.0720 $X2=0.5130 $Y2=0.0720
r10 28 76 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.0720 $X2=0.4840 $Y2=0.0720
r11 32 75 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5130 $Y2=0.0900
r12 73 74 3.78933 $w=1.3e-08 $l=1.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1450 $X2=0.5130 $Y2=0.1612
r13 73 72 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1450 $X2=0.5130 $Y2=0.1217
r14 72 75 7.40378 $w=1.3e-08 $l=3.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1217 $X2=0.5130 $Y2=0.0900
r15 71 74 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1830 $X2=0.5130 $Y2=0.1612
r16 70 71 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5130 $Y2=0.1830
r17 29 33 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2160 $X2=0.5130 $Y2=0.2340
r18 29 70 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2160 $X2=0.5130 $Y2=0.1980
r19 24 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r20 69 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r21 67 66 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r22 23 66 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r23 22 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r24 65 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r25 63 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r26 21 62 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r27 33 61 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.2340 $X2=0.4860 $Y2=0.2340
r28 6 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r29 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3275 $Y2=0.2340
r30 3 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2125 $Y2=0.2340
r31 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1040 $Y2=0.2340
r32 60 61 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r33 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r34 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r35 57 58 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r36 56 57 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3275
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r37 55 56 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3185
+ $Y=0.2340 $X2=0.3275 $Y2=0.2340
r38 54 55 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3185 $Y2=0.2340
r39 53 54 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2605
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r40 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.2340 $X2=0.2605 $Y2=0.2340
r41 51 52 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2215
+ $Y=0.2340 $X2=0.2335 $Y2=0.2340
r42 50 51 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2125
+ $Y=0.2340 $X2=0.2215 $Y2=0.2340
r43 49 50 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.2125 $Y2=0.2340
r44 48 49 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1130
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r45 47 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1040
+ $Y=0.2340 $X2=0.1130 $Y2=0.2340
r46 46 47 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.2340 $X2=0.1040 $Y2=0.2340
r47 27 31 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0540 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r48 27 46 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0855 $Y2=0.2340
r49 31 45 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r50 44 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r51 43 44 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1440 $X2=0.0270 $Y2=0.1980
r52 25 30 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0900 $X2=0.0270 $Y2=0.0720
r53 25 43 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0900 $X2=0.0270 $Y2=0.1440
r54 30 42 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0720 $X2=0.0380 $Y2=0.0720
r55 41 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.0720 $X2=0.0380 $Y2=0.0720
r56 26 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.0720 $X2=0.1080 $Y2=0.0720
r57 26 41 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.0720 $X2=0.0560 $Y2=0.0720
r58 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0720
r59 38 37 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r60 1 37 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r61 34 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.0675 $X2=0.1100 $Y2=0.0675
r62 19 34 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.0980 $Y2=0.0675
r63 35 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r64 4 23 1e-05
r65 2 21 1e-05
.ends


*
.SUBCKT NAND2x2_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@4 N_MM2@4_d N_MM2@4_g N_MM2@4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@4 N_MM3@4_d N_MM3@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@3 N_MM3@3_d N_MM3@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@3 N_MM2@3_d N_MM1@2_g N_MM2@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NAND2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2x2_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2x2_ASAP7_75t_R%noxref_9
cc_1 N_noxref_9_1 N_MM2@2_g 0.001666f
cc_2 N_noxref_9_1 N_NET16_20 0.0361574f
cc_3 N_noxref_9_1 N_Y_20 0.000790826f
x_PM_NAND2x2_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2x2_ASAP7_75t_R%noxref_7
cc_4 N_noxref_7_1 N_MM2_g 0.00166587f
cc_5 N_noxref_7_1 N_NET16_16 0.0362088f
cc_6 N_noxref_7_1 N_Y_19 0.000791236f
x_PM_NAND2x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2x2_ASAP7_75t_R%noxref_10
cc_7 N_noxref_10_1 N_MM2@2_g 0.0091512f
cc_8 N_noxref_10_1 N_NET16_20 0.000638404f
cc_9 N_noxref_10_1 N_Y_29 0.000475855f
cc_10 N_noxref_10_1 N_Y_24 0.00140322f
cc_11 N_noxref_10_1 N_noxref_9_1 0.00193818f
x_PM_NAND2x2_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2x2_ASAP7_75t_R%noxref_8
cc_12 N_noxref_8_1 N_MM2_g 0.00920203f
cc_13 N_noxref_8_1 N_NET16_16 0.000639594f
cc_14 N_noxref_8_1 N_Y_21 0.00183291f
cc_15 N_noxref_8_1 N_noxref_7_1 0.00193398f
x_PM_NAND2x2_ASAP7_75t_R%A VSS A N_MM3_g N_MM3@4_g N_MM3@3_g N_MM0@2_g N_A_7
+ N_A_1 N_A_8 PM_NAND2x2_ASAP7_75t_R%A
cc_16 N_MM0@2_g N_B_12 0.000276878f
cc_17 N_MM0@2_g N_B_1 0.000443022f
cc_18 N_MM0@2_g N_B_2 0.000444752f
cc_19 N_MM0@2_g N_B_10 0.00060935f
cc_20 N_MM0@2_g N_B_19 0.000611778f
cc_21 N_MM0@2_g N_B_14 0.000626726f
cc_22 N_A_7 N_B_12 0.00132999f
cc_23 N_A_1 N_B_12 0.00229684f
cc_24 N_A_7 N_B_21 0.0027246f
cc_25 N_MM3_g N_MM2@4_g 0.00337014f
cc_26 N_MM0@2_g N_MM1@2_g 0.00448849f
x_PM_NAND2x2_ASAP7_75t_R%B VSS B N_MM2_g N_MM2@4_g N_MM1@2_g N_MM2@2_g N_B_12
+ N_B_1 N_B_2 N_B_10 N_B_19 N_B_14 N_B_21 N_B_16 N_B_13 N_B_11 N_B_18 N_B_20
+ N_B_17 N_B_22 N_B_9 N_B_15 PM_NAND2x2_ASAP7_75t_R%B
x_PM_NAND2x2_ASAP7_75t_R%NET16 VSS N_MM2_s N_MM2@4_s N_MM3_d N_MM3@4_d
+ N_MM3@3_d N_MM3@2_d N_MM2@3_s N_MM2@2_s N_NET16_16 N_NET16_21 N_NET16_1
+ N_NET16_5 N_NET16_3 N_NET16_17 N_NET16_20 N_NET16_19 N_NET16_4 N_NET16_2
+ N_NET16_18 PM_NAND2x2_ASAP7_75t_R%NET16
cc_27 N_NET16_16 N_B_16 0.000181707f
cc_28 N_NET16_21 N_B_13 0.000203648f
cc_29 N_NET16_21 N_B_11 0.000207908f
cc_30 N_NET16_1 N_B_1 0.000255426f
cc_31 N_NET16_5 N_B_2 0.000289063f
cc_32 N_NET16_3 N_B_12 0.00112209f
cc_33 N_NET16_17 N_MM2@4_g 0.0335087f
cc_34 N_NET16_20 N_MM2@2_g 0.0340422f
cc_35 N_NET16_19 N_MM1@2_g 0.0336172f
cc_36 N_NET16_21 N_B_18 0.00100858f
cc_37 N_NET16_21 N_B_20 0.00109295f
cc_38 N_NET16_1 N_MM2_g 0.0011198f
cc_39 N_NET16_5 N_MM2@2_g 0.00112071f
cc_40 N_NET16_4 N_B_14 0.00122256f
cc_41 N_NET16_2 N_B_10 0.0012824f
cc_42 N_NET16_4 N_MM1@2_g 0.0014658f
cc_43 N_NET16_2 N_MM2@4_g 0.00148656f
cc_44 N_NET16_20 N_B_2 0.00156308f
cc_45 N_NET16_17 N_B_1 0.00156988f
cc_46 N_NET16_21 N_B_12 0.0110508f
cc_47 N_NET16_16 N_MM2_g 0.0351918f
cc_48 N_NET16_17 N_MM3@3_g 0.000467418f
cc_49 N_NET16_4 N_MM3@3_g 0.000721624f
cc_50 N_NET16_2 N_MM3@3_g 0.000742059f
cc_51 N_NET16_3 N_MM3@3_g 0.0020245f
cc_52 N_NET16_18 N_A_1 0.00376316f
cc_53 N_NET16_19 N_MM0@2_g 0.0330499f
cc_54 N_NET16_17 N_MM3_g 0.0331496f
cc_55 N_NET16_18 N_MM3@4_g 0.0183839f
cc_56 N_NET16_18 N_MM3@3_g 0.0500742f
x_PM_NAND2x2_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM2@4_d N_MM1_d N_MM0_d N_MM0@2_d
+ N_MM1@2_d N_MM2@3_d N_MM2@2_d N_Y_4 N_Y_3 N_Y_2 N_Y_1 N_Y_5 N_Y_6 N_Y_19
+ N_Y_24 N_Y_21 N_Y_26 N_Y_28 N_Y_27 N_Y_25 N_Y_29 N_Y_20 N_Y_23 N_Y_22 N_Y_32
+ N_Y_30 PM_NAND2x2_ASAP7_75t_R%Y
cc_57 N_Y_4 N_MM2@2_g 0.000273173f
cc_58 N_Y_3 N_B_19 0.000160537f
cc_59 N_Y_4 N_MM1@2_g 0.000177622f
cc_60 N_Y_3 N_MM2@4_g 0.000194785f
cc_61 N_Y_2 N_B_17 0.000340913f
cc_62 N_Y_1 N_B_10 0.000424277f
cc_63 N_Y_5 N_B_14 0.000448186f
cc_64 N_Y_2 N_B_1 0.000766819f
cc_65 N_Y_6 N_B_2 0.000882349f
cc_66 N_Y_19 N_MM2@4_g 0.0684021f
cc_67 N_Y_24 N_MM1@2_g 0.0119936f
cc_68 N_Y_21 N_MM2@4_g 0.0328451f
cc_69 N_Y_5 N_MM2@2_g 0.00210326f
cc_70 N_Y_1 N_MM2@4_g 0.00210793f
cc_71 N_Y_26 N_B_10 0.00263182f
cc_72 N_Y_6 N_MM2@2_g 0.00263237f
cc_73 N_Y_28 N_B_14 0.00264566f
cc_74 N_Y_2 N_MM2@4_g 0.00293914f
cc_75 N_Y_27 N_B_17 0.00294386f
cc_76 N_Y_27 N_B_21 0.00389866f
cc_77 N_Y_28 N_B_22 0.00401719f
cc_78 N_Y_26 N_B_16 0.00430423f
cc_79 N_Y_21 N_B_1 0.00461423f
cc_80 N_Y_25 N_B_9 0.00463209f
cc_81 N_Y_24 N_B_2 0.0046579f
cc_82 N_Y_29 N_B_15 0.00489496f
cc_83 N_Y_24 N_MM2@2_g 0.0211752f
cc_84 N_Y_20 N_MM1@2_g 0.0372411f
cc_85 N_Y_19 N_MM2_g 0.0378937f
cc_86 N_Y_20 N_MM2@2_g 0.0697351f
cc_87 N_Y_4 N_MM3@4_g 0.0011028f
cc_88 N_Y_23 N_MM3@4_g 0.00130233f
cc_89 N_Y_4 N_MM0@2_g 0.00256579f
cc_90 N_Y_3 N_MM3@4_g 0.00266629f
cc_91 N_Y_23 N_A_1 0.00514172f
cc_92 N_Y_27 N_A_8 0.00585691f
cc_93 N_Y_23 N_MM3@3_g 0.0193219f
cc_94 N_Y_23 N_MM0@2_g 0.0503415f
cc_95 N_Y_22 N_MM3_g 0.0295259f
cc_96 N_Y_22 N_MM3@4_g 0.0426603f
cc_97 N_Y_1 N_NET16_21 0.000912398f
cc_98 N_Y_5 N_NET16_21 0.000988745f
cc_99 N_Y_26 N_NET16_1 0.000519909f
cc_100 N_Y_28 N_NET16_5 0.000519909f
cc_101 N_Y_20 N_NET16_19 0.000562401f
cc_102 N_Y_19 N_NET16_17 0.00168468f
cc_103 N_Y_32 N_NET16_21 0.000618723f
cc_104 N_Y_30 N_NET16_21 0.000626124f
cc_105 N_Y_19 N_NET16_16 0.000691488f
cc_106 N_Y_20 N_NET16_20 0.0018125f
cc_107 N_Y_29 N_NET16_5 0.000722051f
cc_108 N_Y_25 N_NET16_1 0.000732697f
cc_109 N_Y_5 N_NET16_4 0.00134081f
cc_110 N_Y_1 N_NET16_1 0.00238519f
cc_111 N_Y_26 N_NET16_21 0.00371429f
cc_112 N_Y_28 N_NET16_21 0.00372604f
cc_113 N_Y_1 N_NET16_2 0.0040906f
cc_114 N_Y_5 N_NET16_5 0.00514668f
cc_115 N_Y_4 N_NET16_21 0.00877661f
*END of NAND2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND2xp33_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2xp33_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0317166f
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0208966f
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000842116f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1080 $Y2=0.0540
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00449124f
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0205893f
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%B VSS 4 3 1 6 5
c1 1 VSS 0.000854132f
c2 3 VSS 0.0220841f
c3 4 VSS 0.00434644f
c4 5 VSS 0.0034152f
c5 6 VSS 0.00173642f
r1 6 11 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 5 10 6.11415 $w=1.4371e-08 $l=3.1504e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1345 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 10 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r4 4 11 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1665
r5 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%A VSS 16 3 1 6 5 9
c1 1 VSS 0.00185137f
c2 3 VSS 0.04997f
c3 4 VSS 0.00541831f
c4 5 VSS 0.00508395f
c5 6 VSS 0.00138061f
c6 7 VSS 0.00767673f
c7 8 VSS 0.00108567f
c8 9 VSS 0.00710178f
r1 9 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 7 19 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r5 5 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r6 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 4 18 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 16 6 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r11 16 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r12 12 14 12.3648 $w=1.13e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r13 1 11 3.86521 $w=1.8e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r14 1 12 4.25053 $w=1.32143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r15 3 11 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r16 3 12 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_NAND2xp33_ASAP7_75t_R%Y VSS 18 15 27 28 8 9 1 7 11 2 10
c1 1 VSS 0.0067188f
c2 2 VSS 0.00601127f
c3 7 VSS 0.00303715f
c4 8 VSS 0.00355684f
c5 9 VSS 0.00900671f
c6 10 VSS 0.00397333f
c7 11 VSS 0.00484981f
c8 12 VSS 0.00303428f
c9 13 VSS 0.00363369f
r1 28 26 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2295 $X2=0.1225 $Y2=0.2295
r2 1 26 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2295 $X2=0.1225 $Y2=0.2295
r3 8 1 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2295 $X2=0.1080 $Y2=0.2295
r4 27 8 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2295 $X2=0.0935 $Y2=0.2295
r5 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2295
+ $X2=0.1120 $Y2=0.2340
r6 21 22 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r7 9 13 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2340 $X2=0.1890 $Y2=0.2340
r8 9 22 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r9 13 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r10 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r11 18 19 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1980
r12 18 17 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0720
r13 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0360
r14 11 17 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0720
r15 10 12 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0360 $X2=0.1890 $Y2=0.0360
r16 2 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r17 7 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1600 $Y2=0.0540
r18 15 7 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
.ends


*
.SUBCKT NAND2xp33_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1


*include "NAND2xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2xp33_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2xp33_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM3_g 0.004781f
x_PM_NAND2xp33_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2xp33_ASAP7_75t_R%noxref_8
cc_2 N_noxref_8_1 N_MM3_g 0.00715045f
cc_3 N_noxref_8_1 N_noxref_7_1 0.00202512f
x_PM_NAND2xp33_ASAP7_75t_R%NET16 VSS N_MM3_d N_MM2_s N_NET16_1
+ PM_NAND2xp33_ASAP7_75t_R%NET16
cc_4 N_NET16_1 N_MM3_g 0.0125684f
cc_5 N_NET16_1 N_MM2_g 0.0125438f
x_PM_NAND2xp33_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2xp33_ASAP7_75t_R%noxref_9
cc_6 N_noxref_9_1 N_MM2_g 0.00371889f
cc_7 N_noxref_9_1 N_Y_7 0.0282188f
x_PM_NAND2xp33_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2xp33_ASAP7_75t_R%noxref_10
cc_8 N_noxref_10_1 N_MM2_g 0.00592497f
cc_9 N_noxref_10_1 N_Y_8 0.00138929f
cc_10 N_noxref_10_1 N_noxref_9_1 0.00207849f
x_PM_NAND2xp33_ASAP7_75t_R%B VSS B N_MM2_g N_B_1 N_B_6 N_B_5
+ PM_NAND2xp33_ASAP7_75t_R%B
cc_11 N_B_1 N_A_1 0.00266368f
cc_12 N_B_6 N_A_6 0.000545926f
cc_13 N_B_5 N_A_6 0.000661637f
cc_14 N_B N_A_6 0.00206852f
cc_15 N_MM2_g N_MM3_g 0.0122288f
x_PM_NAND2xp33_ASAP7_75t_R%A VSS A N_MM3_g N_A_1 N_A_6 N_A_5 N_A_9
+ PM_NAND2xp33_ASAP7_75t_R%A
x_PM_NAND2xp33_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM0_d N_MM1_d N_Y_8 N_Y_9 N_Y_1
+ N_Y_7 N_Y_11 N_Y_2 N_Y_10 PM_NAND2xp33_ASAP7_75t_R%Y
cc_16 N_Y_8 N_A_6 0.000222078f
cc_17 N_Y_9 N_A_5 0.000280341f
cc_18 N_Y_1 N_MM3_g 0.000352475f
cc_19 N_Y_9 N_A_9 0.000864317f
cc_20 N_Y_8 N_MM3_g 0.0166268f
cc_21 N_Y_7 N_B_6 0.000375191f
cc_22 N_Y_1 N_MM2_g 0.000482215f
cc_23 N_Y_11 N_B_1 0.000505674f
cc_24 N_Y_7 N_B_1 0.000624555f
cc_25 N_Y_2 N_MM2_g 0.00110197f
cc_26 N_Y_8 N_MM2_g 0.00667028f
cc_27 N_Y_10 N_B_5 0.00261972f
cc_28 N_Y_9 N_B_6 0.00458434f
cc_29 N_Y_11 N_B 0.00628362f
cc_30 N_Y_7 N_MM2_g 0.0345093f
*END of NAND2xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND2xp5_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2xp5_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0419614f
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0321779f
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000930301f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%A VSS 16 3 1 6 9
c1 1 VSS 0.0052945f
c2 3 VSS 0.0714914f
c3 4 VSS 0.00671838f
c4 5 VSS 0.00585688f
c5 6 VSS 0.00169991f
c6 7 VSS 0.00803618f
c7 8 VSS 0.00134786f
c8 9 VSS 0.00710778f
r1 9 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 7 19 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r5 5 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r6 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 4 18 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 16 6 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r11 16 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r12 12 14 12.3648 $w=1.13e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r13 1 11 3.86521 $w=1.8e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r14 1 12 4.25053 $w=1.32143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r15 3 11 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r16 3 12 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00489003f
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0316045f
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%B VSS 12 3 1 6 5 4
c1 1 VSS 0.00131948f
c2 3 VSS 0.0328078f
c3 4 VSS 0.0057786f
c4 5 VSS 0.00423941f
c5 6 VSS 0.00219366f
r1 6 13 5.17411 $w=1.46514e-08 $l=2.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1707
r2 5 10 6.11415 $w=1.4371e-08 $l=3.1504e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1345 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 12 13 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1520 $X2=0.1350 $Y2=0.1707
r4 12 11 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1520 $X2=0.1350 $Y2=0.1477
r5 4 10 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r6 4 11 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1477
r7 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r8 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NAND2xp5_ASAP7_75t_R%Y VSS 19 15 30 31 8 1 9 7 2 10 11
c1 1 VSS 0.00887324f
c2 2 VSS 0.00638375f
c3 7 VSS 0.00286293f
c4 8 VSS 0.00407343f
c5 9 VSS 0.00905067f
c6 10 VSS 0.00387141f
c7 11 VSS 0.00428447f
c8 12 VSS 0.00296044f
c9 13 VSS 0.00345922f
r1 31 29 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 1 29 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 8 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 30 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1120 $Y2=0.2340
r6 23 24 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r7 9 13 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2340 $X2=0.1890 $Y2=0.2340
r8 9 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r9 13 22 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r10 21 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r11 20 21 14.3995 $w=1.3e-08 $l=6.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1362 $X2=0.1890 $Y2=0.1980
r12 19 20 12.4174 $w=1.3e-08 $l=5.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0830 $X2=0.1890 $Y2=0.1362
r13 19 18 0.291487 $w=1.3e-08 $l=1.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0830 $X2=0.1890 $Y2=0.0817
r14 17 18 2.2736 $w=1.3e-08 $l=9.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0720 $X2=0.1890 $Y2=0.0817
r15 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0360
r16 11 17 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0720
r17 10 12 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0360 $X2=0.1890 $Y2=0.0360
r18 2 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r19 7 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r20 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
.ends


*
.SUBCKT NAND2xp5_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND2xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2xp5_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2xp5_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM3_g 0.00255734f
x_PM_NAND2xp5_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2xp5_ASAP7_75t_R%noxref_8
cc_2 N_noxref_8_1 N_MM3_g 0.00463163f
cc_3 N_noxref_8_1 N_noxref_7_1 0.00186189f
x_PM_NAND2xp5_ASAP7_75t_R%NET16 VSS N_MM3_d N_MM2_s N_NET16_1
+ PM_NAND2xp5_ASAP7_75t_R%NET16
cc_4 N_NET16_1 N_MM3_g 0.0173744f
cc_5 N_NET16_1 N_MM2_g 0.0174044f
x_PM_NAND2xp5_ASAP7_75t_R%A VSS A N_MM3_g N_A_1 N_A_6 N_A_9
+ PM_NAND2xp5_ASAP7_75t_R%A
x_PM_NAND2xp5_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2xp5_ASAP7_75t_R%noxref_9
cc_6 N_noxref_9_1 N_MM2_g 0.00162212f
cc_7 N_noxref_9_1 N_Y_7 0.0379425f
x_PM_NAND2xp5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2xp5_ASAP7_75t_R%noxref_10
cc_8 N_noxref_10_1 N_MM2_g 0.00349817f
cc_9 N_noxref_10_1 N_Y_8 0.00156052f
cc_10 N_noxref_10_1 N_noxref_9_1 0.00189393f
x_PM_NAND2xp5_ASAP7_75t_R%B VSS B N_MM2_g N_B_1 N_B_6 N_B_5 N_B_4
+ PM_NAND2xp5_ASAP7_75t_R%B
cc_11 N_B_1 N_A_1 0.00216478f
cc_12 N_B_6 N_A_6 0.000476648f
cc_13 N_B_5 N_A_6 0.000614698f
cc_14 N_B_4 N_A_6 0.00192472f
cc_15 N_MM2_g N_MM3_g 0.00854719f
x_PM_NAND2xp5_ASAP7_75t_R%Y VSS Y N_MM2_d N_MM0_d N_MM1_d N_Y_8 N_Y_1 N_Y_9
+ N_Y_7 N_Y_2 N_Y_10 N_Y_11 PM_NAND2xp5_ASAP7_75t_R%Y
cc_16 N_Y_8 N_A_1 0.000364732f
cc_17 N_Y_1 N_MM3_g 0.000574459f
cc_18 N_Y_9 N_A_9 0.000876636f
cc_19 N_Y_8 N_MM3_g 0.0267792f
cc_20 N_Y_7 N_B_1 0.00184876f
cc_21 N_Y_1 N_MM2_g 0.000910862f
cc_22 N_Y_2 N_MM2_g 0.00183973f
cc_23 N_Y_10 N_B_5 0.00257866f
cc_24 N_Y_8 N_MM2_g 0.0109762f
cc_25 N_Y_9 N_B_6 0.0044647f
cc_26 N_Y_11 N_B_4 0.0063883f
cc_27 N_Y_7 N_MM2_g 0.050227f
*END of NAND2xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND2xp67_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND2xp67_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND2xp67_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND2xp67_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0318832f
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00503173f
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00485072f
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00509874f
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%B VSS 21 3 4 1 5 6
c1 1 VSS 0.00653487f
c2 3 VSS 0.0342394f
c3 4 VSS 0.035628f
c4 5 VSS 0.00341501f
c5 6 VSS 0.0036704f
r1 6 22 4.70773 $w=1.47822e-08 $l=2.53e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1980 $X2=0.2430 $Y2=0.1727
r2 21 22 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1560 $X2=0.2430 $Y2=0.1727
r3 21 20 1.45744 $w=1.3e-08 $l=6.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1560 $X2=0.2430 $Y2=0.1497
r4 19 20 1.45744 $w=1.3e-08 $l=6.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1435 $X2=0.2430 $Y2=0.1497
r5 17 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1345 $X2=0.2430 $Y2=0.1435
r6 5 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1255 $X2=0.2430 $Y2=0.1345
r7 4 14 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1340
r8 14 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1340
+ $X2=0.2430 $Y2=0.1345
r9 13 14 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1340 $X2=0.2430 $Y2=0.1340
r10 11 13 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1340 $X2=0.2335 $Y2=0.1340
r11 10 11 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1340 $X2=0.2305 $Y2=0.1340
r12 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1340 $X2=0.2160 $Y2=0.1340
r13 3 1 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1340
r14 1 8 3.05464 $w=2.15326e-08 $l=1.08e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1340 $X2=0.1782 $Y2=0.1340
r15 1 9 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1340 $X2=0.2015 $Y2=0.1340
r16 3 8 0.757708 $w=2.1223e-07 $l=1.08462e-08 $layer=LIG $thickness=5.54419e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1782 $Y2=0.1340
r17 3 9 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1340
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%Y VSS 27 17 20 41 43 9 1 10 2 12 8 11 13 14
c1 1 VSS 0.013227f
c2 2 VSS 0.00291928f
c3 8 VSS 0.00213661f
c4 9 VSS 0.00295848f
c5 10 VSS 0.00285113f
c6 11 VSS 0.0148391f
c7 12 VSS 0.000843198f
c8 13 VSS 0.00254993f
c9 14 VSS 0.000773281f
c10 15 VSS 0.00302279f
r1 9 38 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1060 $Y2=0.2160
r2 43 9 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r3 41 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 10 40 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 38 39 3.74659 $w=5.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1080 $Y=0.2160 $X2=0.1330 $Y2=0.2160
r6 37 39 2.24795 $w=5.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1480 $Y=0.2160 $X2=0.1330 $Y2=0.2160
r7 1 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r8 1 37 2.09809 $w=5.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08 $X=0.1620
+ $Y=0.2160 $X2=0.1480 $Y2=0.2160
r9 35 36 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1865 $Y2=0.2340
r10 33 36 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2085
+ $Y=0.2340 $X2=0.1865 $Y2=0.2340
r11 32 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.2340 $X2=0.2085 $Y2=0.2340
r12 11 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2970 $Y2=0.2340
r13 11 32 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2335 $Y2=0.2340
r14 15 31 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2970 $Y2=0.2160
r15 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2970 $Y2=0.2160
r16 29 30 11.7178 $w=1.3e-08 $l=5.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1477 $X2=0.2970 $Y2=0.1980
r17 28 29 9.67738 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1062 $X2=0.2970 $Y2=0.1477
r18 27 28 0.116595 $w=1.3e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1057 $X2=0.2970 $Y2=0.1062
r19 27 13 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1057 $X2=0.2970 $Y2=0.0932
r20 13 14 3.30617 $w=1.71506e-08 $l=2.12e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0932 $X2=0.2970 $Y2=0.0720
r21 14 26 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0720 $X2=0.2860 $Y2=0.0720
r22 25 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2680
+ $Y=0.0720 $X2=0.2860 $Y2=0.0720
r23 24 25 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0720 $X2=0.2680 $Y2=0.0720
r24 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r25 22 23 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2200
+ $Y=0.0720 $X2=0.2295 $Y2=0.0720
r26 21 22 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2110
+ $Y=0.0720 $X2=0.2200 $Y2=0.0720
r27 12 21 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0720 $X2=0.2110 $Y2=0.0720
r28 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2200 $Y2=0.0720
r29 20 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r30 18 19 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r31 2 18 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0540 $X2=0.2260 $Y2=0.0540
r32 8 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2140 $Y2=0.0540
r33 17 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r34 1 10 1e-05
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%NET15 VSS 15 27 30 32 1 2 10 13 11 3 12
c1 1 VSS 0.00759319f
c2 2 VSS 0.00645428f
c3 3 VSS 0.00483185f
c4 10 VSS 0.00322869f
c5 11 VSS 0.0029474f
c6 12 VSS 0.00222109f
c7 13 VSS 0.0224072f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0540 $X2=0.2680 $Y2=0.0540
r2 32 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2555 $Y2=0.0540
r3 30 29 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r4 2 29 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r5 26 2 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.0540 $X2=0.1640 $Y2=0.0540
r6 11 26 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1520 $Y2=0.0540
r7 27 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r8 3 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r9 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r10 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r11 22 23 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1865
+ $Y=0.0360 $X2=0.2315 $Y2=0.0360
r12 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1865 $Y2=0.0360
r13 20 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r14 19 20 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1505 $Y2=0.0360
r15 18 19 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r16 17 18 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.0360 $X2=0.0790 $Y2=0.0360
r17 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.0360 $X2=0.0590 $Y2=0.0360
r18 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0500 $Y2=0.0360
r19 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0500 $Y2=0.0360
r20 15 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r21 10 14 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r22 1 10 1e-05
.ends

.subckt PM_NAND2xp67_ASAP7_75t_R%A VSS 22 3 4 8 1
c1 1 VSS 0.00323685f
c2 3 VSS 0.0593146f
c3 4 VSS 0.0318144f
c4 5 VSS 0.00364932f
c5 6 VSS 0.00845178f
c6 7 VSS 0.00298268f
c7 8 VSS 0.00373893f
c8 9 VSS 0.00183577f
c9 10 VSS 0.00882485f
r1 10 27 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 8 25 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0720 $X2=0.0270 $Y2=0.0935
r3 26 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 6 9 6.28176 $w=1.44063e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1660 $X2=0.0270 $Y2=0.1340
r5 6 26 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1660 $X2=0.0270 $Y2=0.1980
r6 5 9 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1155 $X2=0.0270 $Y2=0.1340
r7 5 25 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1155 $X2=0.0270 $Y2=0.0935
r8 9 24 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1340 $X2=0.0455 $Y2=0.1340
r9 4 20 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1340
r10 22 7 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0635 $Y2=0.1340
r11 7 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1340 $X2=0.0455 $Y2=0.1340
r12 18 20 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1340 $X2=0.1350 $Y2=0.1340
r13 17 18 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1340 $X2=0.1225 $Y2=0.1340
r14 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1340 $X2=0.1080 $Y2=0.1340
r15 13 16 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1340 $X2=0.0935 $Y2=0.1340
r16 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0905 $Y2=0.1340
r17 22 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1340
+ $X2=0.0810 $Y2=0.1340
r18 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1340 $X2=0.0810 $Y2=0.1340
r19 1 14 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0715 $Y=0.1340 $X2=0.0685 $Y2=0.1340
r20 3 12 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1340
r21 3 14 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1340
r22 3 16 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1340
.ends


*
.SUBCKT NAND2xp67_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4@2 N_MM4@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3@2 N_MM3@2_d N_MM3@2_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND2xp67_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND2xp67_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND2xp67_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NAND2xp67_ASAP7_75t_R%noxref_8
cc_1 N_noxref_8_1 N_MM4_g 0.00469376f
cc_2 N_noxref_8_1 N_noxref_7_1 0.0020318f
x_PM_NAND2xp67_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NAND2xp67_ASAP7_75t_R%noxref_7
cc_3 N_noxref_7_1 N_MM4_g 0.00460377f
cc_4 N_noxref_7_1 N_NET15_10 0.0269635f
x_PM_NAND2xp67_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND2xp67_ASAP7_75t_R%noxref_9
cc_5 N_noxref_9_1 N_MM3@2_g 0.00376459f
cc_6 N_noxref_9_1 N_NET15_12 0.0268736f
cc_7 N_noxref_9_1 N_Y_8 0.000929665f
x_PM_NAND2xp67_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND2xp67_ASAP7_75t_R%noxref_10
cc_8 N_noxref_10_1 N_MM3@2_g 0.00952812f
cc_9 N_noxref_10_1 N_NET15_12 0.00018594f
cc_10 N_noxref_10_1 N_Y_13 0.00133623f
cc_11 N_noxref_10_1 N_noxref_9_1 0.00210324f
x_PM_NAND2xp67_ASAP7_75t_R%B VSS B N_MM3_g N_MM3@2_g N_B_1 N_B_5 N_B_6
+ PM_NAND2xp67_ASAP7_75t_R%B
cc_12 N_B_1 N_MM4@2_g 0.00191989f
cc_13 N_MM3_g N_MM4@2_g 0.00822792f
x_PM_NAND2xp67_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM3@2_d N_MM5_d N_MM2_d N_Y_9
+ N_Y_1 N_Y_10 N_Y_2 N_Y_12 N_Y_8 N_Y_11 N_Y_13 N_Y_14
+ PM_NAND2xp67_ASAP7_75t_R%Y
cc_14 N_Y_9 N_MM4_g 0.0228518f
cc_15 N_Y_9 N_A_1 0.00121929f
cc_16 N_Y_1 N_MM4@2_g 0.00245551f
cc_17 N_Y_9 N_MM4@2_g 0.0147224f
cc_18 N_Y_10 N_MM4@2_g 0.0418816f
cc_19 N_Y_1 N_MM3_g 0.000696668f
cc_20 N_Y_2 N_MM3@2_g 0.000867708f
cc_21 N_Y_12 N_B_5 0.00142387f
cc_22 N_Y_8 N_B_1 0.00169068f
cc_23 N_Y_10 N_MM3_g 0.0108779f
cc_24 N_Y_11 N_B_6 0.00490886f
cc_25 N_Y_13 N_B_5 0.00585071f
cc_26 N_Y_8 N_MM3@2_g 0.0356421f
cc_27 N_Y_8 N_MM3_g 0.0298212f
cc_28 N_Y_12 N_NET15_12 0.000516913f
cc_29 N_Y_12 N_NET15_3 0.000559404f
cc_30 N_Y_14 N_NET15_13 0.000592603f
cc_31 N_Y_2 N_NET15_13 0.000773427f
cc_32 N_Y_8 N_NET15_12 0.000834817f
cc_33 N_Y_2 N_NET15_2 0.00106223f
cc_34 N_Y_2 N_NET15_3 0.003858f
cc_35 N_Y_12 N_NET15_13 0.00968801f
x_PM_NAND2xp67_ASAP7_75t_R%NET15 VSS N_MM4_d N_MM4@2_d N_MM3_s N_MM3@2_s
+ N_NET15_1 N_NET15_2 N_NET15_10 N_NET15_13 N_NET15_11 N_NET15_3 N_NET15_12
+ PM_NAND2xp67_ASAP7_75t_R%NET15
cc_36 N_NET15_1 N_MM4@2_g 0.0004123f
cc_37 N_NET15_2 N_MM4@2_g 0.000528717f
cc_38 N_NET15_1 N_A_8 0.00053619f
cc_39 N_NET15_10 N_A_1 0.000981742f
cc_40 N_NET15_1 N_MM4_g 0.00127053f
cc_41 N_NET15_13 N_MM4@2_g 0.00195214f
cc_42 N_NET15_13 N_A_8 0.00210551f
cc_43 N_NET15_10 N_MM4_g 0.0243646f
cc_44 N_NET15_11 N_MM4@2_g 0.0258952f
cc_45 N_NET15_2 N_MM3_g 0.000528462f
cc_46 N_NET15_3 N_MM3@2_g 0.000556941f
cc_47 N_NET15_12 N_B_1 0.000667438f
cc_48 N_NET15_12 N_MM3@2_g 0.0242627f
cc_49 N_NET15_11 N_MM3_g 0.0257768f
x_PM_NAND2xp67_ASAP7_75t_R%A VSS A N_MM4_g N_MM4@2_g N_A_8 N_A_1
+ PM_NAND2xp67_ASAP7_75t_R%A
*END of NAND2xp67_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND3x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND3x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND3x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND3x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00588155f
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0423497f
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%NET21 VSS 16 17 32 33 36 37 10 1 11 12 3 13 2
c1 1 VSS 0.00980755f
c2 2 VSS 0.0063484f
c3 3 VSS 0.00318603f
c4 10 VSS 0.00447361f
c5 11 VSS 0.00342389f
c6 12 VSS 0.00210418f
c7 13 VSS 0.0131705f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r2 3 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r4 36 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r5 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r6 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r8 32 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r9 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0720
r10 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r11 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0720 $X2=0.3240 $Y2=0.0720
r12 26 27 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2810
+ $Y=0.0720 $X2=0.3105 $Y2=0.0720
r13 25 26 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2510
+ $Y=0.0720 $X2=0.2810 $Y2=0.0720
r14 24 25 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2445
+ $Y=0.0720 $X2=0.2510 $Y2=0.0720
r15 23 24 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2340
+ $Y=0.0720 $X2=0.2445 $Y2=0.0720
r16 22 23 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.2340 $Y2=0.0720
r17 21 22 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r18 20 21 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0720 $X2=0.2045 $Y2=0.0720
r19 19 20 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.0720 $X2=0.1890 $Y2=0.0720
r20 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0720 $X2=0.1465 $Y2=0.0720
r21 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0720 $X2=0.1080 $Y2=0.0720
r22 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0720
r23 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r24 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r25 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r26 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00468072f
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00535479f
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%C VSS 24 3 4 5 6 1
c1 1 VSS 0.0211904f
c2 3 VSS 0.0492408f
c3 4 VSS 0.0858723f
c4 5 VSS 0.084136f
c5 6 VSS 0.0095768f
r1 5 21 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 4 15 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 24 6 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0700 $Y2=0.1170
r4 19 21 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 18 19 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r6 16 18 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r7 15 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r8 13 15 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r9 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r10 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r11 1 7 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1350 $X2=0.0850 $Y2=0.1350
r12 1 8 3.76121 $w=1.74231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0750 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r13 24 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1350
r14 3 7 2.2201 $w=1.49375e-07 $l=4e-09 $layer=LIG $thickness=5.3e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0850 $Y2=0.1350
r15 3 8 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r16 3 11 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%A VSS 8 3 4 5 1 10 6 9 7
c1 1 VSS 0.0095498f
c2 3 VSS 0.0464287f
c3 4 VSS 0.00901001f
c4 5 VSS 0.00990761f
c5 6 VSS 0.00483905f
c6 7 VSS 0.00509465f
c7 8 VSS 0.00420471f
c8 9 VSS 0.00397415f
c9 10 VSS 0.00411086f
r1 7 10 6.04615 $w=1.43636e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4260 $Y=0.1890 $X2=0.4590 $Y2=0.1890
r2 6 9 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.1170 $X2=0.4590 $Y2=0.1170
r3 10 25 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1890 $X2=0.4590 $Y2=0.1620
r4 5 23 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 8 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1620
r6 8 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r7 8 9 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1170
r8 4 17 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r9 21 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r10 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r11 18 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r12 17 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r13 15 17 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r14 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r15 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r16 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r17 1 12 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r18 1 13 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r19 3 12 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r20 3 13 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%NET22 VSS 15 18 29 32 35 36 1 10 11 12 3 2 13
c1 1 VSS 0.00451955f
c2 2 VSS 0.00448122f
c3 3 VSS 0.00450066f
c4 10 VSS 0.00210642f
c5 11 VSS 0.0020885f
c6 12 VSS 0.00205273f
c7 13 VSS 0.0204204f
r1 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r2 3 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r4 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r5 32 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r6 2 31 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r7 28 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3680 $Y=0.0675 $X2=0.3800 $Y2=0.0675
r8 11 28 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3680 $Y2=0.0675
r9 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r10 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r11 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r12 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r13 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4090
+ $Y=0.0360 $X2=0.4475 $Y2=0.0360
r14 23 24 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3935
+ $Y=0.0360 $X2=0.4090 $Y2=0.0360
r15 22 23 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3935 $Y2=0.0360
r16 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r17 20 21 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.0360 $X2=0.3535 $Y2=0.0360
r18 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3085 $Y2=0.0360
r19 13 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r20 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r21 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r22 16 17 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r23 1 16 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.0675 $X2=0.2800 $Y2=0.0675
r24 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r25 15 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%B VSS 8 3 4 5 9 1 7 6 10
c1 1 VSS 0.0149863f
c2 3 VSS 0.046199f
c3 4 VSS 0.0482661f
c4 5 VSS 0.0484312f
c5 6 VSS 0.00585412f
c6 7 VSS 0.00455587f
c7 8 VSS 0.00488634f
c8 9 VSS 0.00407463f
c9 10 VSS 0.0047079f
r1 6 10 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2670
+ $Y=0.1890 $X2=0.2970 $Y2=0.1890
r2 7 9 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2670
+ $Y=0.1170 $X2=0.2970 $Y2=0.1170
r3 10 25 4.64701 $w=1.62667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1890 $X2=0.2970 $Y2=0.1620
r4 5 23 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 8 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1620
r6 8 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r7 8 9 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1170
r8 4 17 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 21 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r10 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r11 18 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r12 17 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r13 15 17 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r14 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r15 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r16 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r17 1 12 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r18 1 13 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r19 3 12 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r20 3 13 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NAND3x1_ASAP7_75t_R%Y VSS 34 23 26 38 50 53 54 1 15 17 2 4 3 19 16
+ 18 14 13
c1 1 VSS 0.0113224f
c2 2 VSS 0.00288853f
c3 3 VSS 0.00760083f
c4 4 VSS 0.0040953f
c5 13 VSS 0.002152f
c6 14 VSS 0.00232659f
c7 15 VSS 0.0047664f
c8 16 VSS 0.00347008f
c9 17 VSS 0.0350005f
c10 18 VSS 0.00210798f
c11 19 VSS 0.00272901f
c12 20 VSS 0.00108931f
c13 21 VSS 0.00258317f
r1 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 1 52 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 15 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 54 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 16 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r6 50 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r7 1 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r8 3 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r9 47 48 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2340 $Y2=0.2340
r10 45 48 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2745
+ $Y=0.2340 $X2=0.2340 $Y2=0.2340
r11 44 45 11.0765 $w=1.3e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.2340 $X2=0.2745 $Y2=0.2340
r12 43 44 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3690
+ $Y=0.2340 $X2=0.3220 $Y2=0.2340
r13 42 43 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4010
+ $Y=0.2340 $X2=0.3690 $Y2=0.2340
r14 40 41 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4545 $Y2=0.2340
r15 39 40 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4125
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r16 39 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4125
+ $Y=0.2340 $X2=0.4010 $Y2=0.2340
r17 17 21 10.9431 $w=1.38333e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.2340 $X2=0.5670 $Y2=0.2340
r18 17 41 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.4545 $Y2=0.2340
r19 21 36 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.2340 $X2=0.5670 $Y2=0.2115
r20 14 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5380 $Y2=0.0675
r21 38 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r22 35 36 9.50248 $w=1.3e-08 $l=4.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1707 $X2=0.5670 $Y2=0.2115
r23 34 35 6.47102 $w=1.3e-08 $l=2.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1430 $X2=0.5670 $Y2=0.1707
r24 34 33 4.13912 $w=1.3e-08 $l=1.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1430 $X2=0.5670 $Y2=0.1252
r25 19 20 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0945 $X2=0.5670 $Y2=0.0720
r26 19 33 7.17059 $w=1.3e-08 $l=3.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0945 $X2=0.5670 $Y2=0.1252
r27 4 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0720
r28 20 32 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0720 $X2=0.5535 $Y2=0.0720
r29 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0720 $X2=0.5535 $Y2=0.0720
r30 30 31 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5155
+ $Y=0.0720 $X2=0.5400 $Y2=0.0720
r31 29 30 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.0720 $X2=0.5155 $Y2=0.0720
r32 28 29 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4545
+ $Y=0.0720 $X2=0.4840 $Y2=0.0720
r33 27 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0720 $X2=0.4545 $Y2=0.0720
r34 18 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0720 $X2=0.4320 $Y2=0.0720
r35 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0720
r36 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r37 24 25 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r38 2 24 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.0675 $X2=0.4420 $Y2=0.0675
r39 13 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r40 23 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
.ends


*
.SUBCKT NAND3x1_ASAP7_75t_R VSS VDD C B A Y
*
* VSS VSS
* VDD VDD
* C C
* B B
* A A
* Y Y
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@3 N_MM2@3_d N_MM2@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM4_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@3 N_MM1@3_d N_MM1@3_g N_MM1@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 N_MM0@3_d N_MM0@3_g N_MM0@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g N_MM0@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NAND3x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND3x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND3x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND3x1_ASAP7_75t_R%noxref_10
cc_1 N_noxref_10_1 N_MM2_g 0.0102683f
cc_2 N_noxref_10_1 N_noxref_9_1 0.00195037f
x_PM_NAND3x1_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND3x1_ASAP7_75t_R%noxref_9
cc_3 N_noxref_9_1 N_MM2_g 0.00200579f
x_PM_NAND3x1_ASAP7_75t_R%NET21 VSS N_MM2_d N_MM2@3_d N_MM2@2_d N_MM1_s
+ N_MM1@3_s N_MM1@2_s N_NET21_10 N_NET21_1 N_NET21_11 N_NET21_12 N_NET21_3
+ N_NET21_13 N_NET21_2 PM_NAND3x1_ASAP7_75t_R%NET21
cc_4 N_NET21_10 N_C_6 0.000973667f
cc_5 N_NET21_10 N_C_1 0.00447271f
cc_6 N_NET21_1 N_MM2@3_g 0.00177553f
cc_7 N_NET21_11 N_MM2@2_g 0.0325733f
cc_8 N_NET21_10 N_MM2_g 0.0181248f
cc_9 N_NET21_10 N_MM2@3_g 0.0497341f
cc_10 N_NET21_12 N_B_9 0.00107334f
cc_11 N_NET21_3 N_MM1@2_g 0.00182481f
cc_12 N_NET21_12 N_B_1 0.00320089f
cc_13 N_NET21_13 N_B_7 0.00439948f
cc_14 N_NET21_11 N_MM4_g 0.0326226f
cc_15 N_NET21_12 N_MM1@3_g 0.01814f
cc_16 N_NET21_12 N_MM1@2_g 0.0505691f
x_PM_NAND3x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NAND3x1_ASAP7_75t_R%noxref_12
cc_17 N_noxref_12_1 N_MM0@2_g 0.00942774f
cc_18 N_noxref_12_1 N_Y_14 0.00216859f
cc_19 N_noxref_12_1 N_noxref_11_1 0.00193687f
x_PM_NAND3x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NAND3x1_ASAP7_75t_R%noxref_11
cc_20 N_noxref_11_1 N_MM0@2_g 0.00164944f
cc_21 N_noxref_11_1 N_Y_14 0.03738f
x_PM_NAND3x1_ASAP7_75t_R%C VSS C N_MM2_g N_MM2@3_g N_MM2@2_g N_C_6 N_C_1
+ PM_NAND3x1_ASAP7_75t_R%C
x_PM_NAND3x1_ASAP7_75t_R%A VSS A N_MM3_g N_MM0@3_g N_MM0@2_g N_A_1 N_A_10 N_A_6
+ N_A_9 N_A_7 PM_NAND3x1_ASAP7_75t_R%A
cc_22 N_MM3_g N_MM1@2_g 0.00550386f
x_PM_NAND3x1_ASAP7_75t_R%NET22 VSS N_MM1_d N_MM1@3_d N_MM1@2_d N_MM0_s
+ N_MM0@3_s N_MM0@2_s N_NET22_1 N_NET22_10 N_NET22_11 N_NET22_12 N_NET22_3
+ N_NET22_2 N_NET22_13 PM_NAND3x1_ASAP7_75t_R%NET22
cc_23 N_NET22_1 N_MM1@3_g 0.00196472f
cc_24 N_NET22_10 N_B_1 0.00288571f
cc_25 N_NET22_11 N_MM1@2_g 0.0325775f
cc_26 N_NET22_10 N_MM4_g 0.0180227f
cc_27 N_NET22_10 N_MM1@3_g 0.0502689f
cc_28 N_NET22_12 N_MM3_g 0.000920729f
cc_29 N_NET22_3 N_MM0@2_g 0.00176066f
cc_30 N_NET22_12 N_A_1 0.00271512f
cc_31 N_NET22_11 N_MM3_g 0.0327059f
cc_32 N_NET22_12 N_MM0@3_g 0.018107f
cc_33 N_NET22_12 N_MM0@2_g 0.0498933f
cc_34 N_NET22_11 N_NET21_13 0.0011066f
cc_35 N_NET22_10 N_NET21_12 0.0011158f
cc_36 N_NET22_1 N_NET21_2 0.00123326f
cc_37 N_NET22_1 N_NET21_3 0.00301238f
cc_38 N_NET22_2 N_NET21_3 0.00416378f
cc_39 N_NET22_13 N_NET21_13 0.0117862f
x_PM_NAND3x1_ASAP7_75t_R%B VSS B N_MM4_g N_MM1@3_g N_MM1@2_g N_B_9 N_B_1 N_B_7
+ N_B_6 N_B_10 PM_NAND3x1_ASAP7_75t_R%B
cc_40 N_MM4_g N_MM2@2_g 0.00490617f
x_PM_NAND3x1_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM0@3_d N_MM0@2_d N_MM3_d N_MM4_d
+ N_MM5_d N_Y_1 N_Y_15 N_Y_17 N_Y_2 N_Y_4 N_Y_3 N_Y_19 N_Y_16 N_Y_18 N_Y_14
+ N_Y_13 PM_NAND3x1_ASAP7_75t_R%Y
cc_41 N_Y_1 N_MM2@2_g 0.000803783f
cc_42 N_Y_15 N_C_1 0.000915891f
cc_43 N_Y_15 N_MM2@2_g 0.0343346f
cc_44 N_Y_15 N_B_1 0.000983479f
cc_45 N_Y_1 N_MM4_g 0.00114261f
cc_46 N_Y_17 N_B_6 0.00185745f
cc_47 N_Y_17 N_B_10 0.00378389f
cc_48 N_Y_15 N_MM4_g 0.0353115f
cc_49 N_Y_2 N_MM0@3_g 0.00241457f
cc_50 N_Y_4 N_MM0@2_g 0.000875919f
cc_51 N_Y_3 N_A 0.00100495f
cc_52 N_Y_19 N_A_1 0.00119459f
cc_53 N_Y_16 N_MM3_g 0.0119303f
cc_54 N_Y_17 N_A_10 0.00129324f
cc_55 N_Y_18 N_A_6 0.00173767f
cc_56 N_Y_3 N_MM0@3_g 0.00308861f
cc_57 N_Y_18 N_A_9 0.0034473f
cc_58 N_Y_17 N_A_7 0.00532738f
cc_59 N_Y_16 N_A_1 0.00601792f
cc_60 N_Y_14 N_MM0@2_g 0.0347333f
cc_61 N_Y_16 N_MM0@3_g 0.0211654f
cc_62 N_Y_13 N_MM3_g 0.0372387f
cc_63 N_Y_13 N_MM0@3_g 0.0699354f
cc_64 N_Y_14 N_NET22_13 0.000552902f
cc_65 N_Y_13 N_NET22_13 0.000560096f
cc_66 N_Y_2 N_NET22_13 0.00069004f
cc_67 N_Y_13 N_NET22_12 0.00111006f
cc_68 N_Y_14 N_NET22_12 0.00111936f
cc_69 N_Y_2 N_NET22_2 0.00134233f
cc_70 N_Y_2 N_NET22_3 0.00279336f
cc_71 N_Y_4 N_NET22_3 0.00441352f
cc_72 N_Y_18 N_NET22_13 0.0101712f
*END of NAND3x1_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND3x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND3x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND3x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND3x2_ASAP7_75t_R%NET21 VSS 28 29 53 54 57 58 61 62 65 66 69 70 24
+ 20 4 19 5 2 1 6 25 23 22 3 21
c1 1 VSS 0.00310225f
c2 2 VSS 0.00609197f
c3 3 VSS 0.00953536f
c4 4 VSS 0.00954848f
c5 5 VSS 0.00617838f
c6 6 VSS 0.00335351f
c7 19 VSS 0.0021165f
c8 20 VSS 0.00338633f
c9 21 VSS 0.00437076f
c10 22 VSS 0.00436397f
c11 23 VSS 0.00336268f
c12 24 VSS 0.00211297f
c13 25 VSS 0.0333981f
r1 70 68 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.0675 $X2=0.8245 $Y2=0.0675
r2 6 68 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.0675 $X2=0.8245 $Y2=0.0675
r3 24 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8100 $Y2=0.0675
r4 69 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r5 66 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r6 5 64 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r7 23 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r8 65 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r9 62 60 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r10 1 60 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r11 19 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r12 61 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r13 58 56 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r14 2 56 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r15 20 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r16 57 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r17 54 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r18 3 52 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r19 21 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r20 53 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r21 6 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0675
+ $X2=0.8100 $Y2=0.0720
r22 5 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0675
+ $X2=0.7020 $Y2=0.0720
r23 1 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0720
r24 2 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0720
r25 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0720
r26 48 49 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7720
+ $Y=0.0720 $X2=0.8100 $Y2=0.0720
r27 47 48 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.0720 $X2=0.7720 $Y2=0.0720
r28 46 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7335
+ $Y=0.0720 $X2=0.7425 $Y2=0.0720
r29 45 46 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7180
+ $Y=0.0720 $X2=0.7335 $Y2=0.0720
r30 44 45 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0720 $X2=0.7180 $Y2=0.0720
r31 43 44 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6775
+ $Y=0.0720 $X2=0.7020 $Y2=0.0720
r32 42 43 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6325
+ $Y=0.0720 $X2=0.6775 $Y2=0.0720
r33 41 42 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0720 $X2=0.6325 $Y2=0.0720
r34 40 41 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5750
+ $Y=0.0720 $X2=0.5940 $Y2=0.0720
r35 38 39 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0720 $X2=0.3085 $Y2=0.0720
r36 36 39 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.0720 $X2=0.3085 $Y2=0.0720
r37 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0720 $X2=0.4025 $Y2=0.0720
r38 33 34 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3625
+ $Y=0.0720 $X2=0.3780 $Y2=0.0720
r39 33 36 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3625
+ $Y=0.0720 $X2=0.3470 $Y2=0.0720
r40 31 32 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0720 $X2=0.5210 $Y2=0.0720
r41 30 31 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0720 $X2=0.4860 $Y2=0.0720
r42 30 35 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.0720 $X2=0.4025 $Y2=0.0720
r43 25 32 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.0720 $X2=0.5210 $Y2=0.0720
r44 25 40 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.0720 $X2=0.5750 $Y2=0.0720
r45 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0720
r46 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r47 4 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r48 22 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r49 29 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00534627f
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00468242f
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00468447f
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%NET22__2 VSS 16 17 29 32 34 37 10 2 1 11 12 3 13
c1 1 VSS 0.00434496f
c2 2 VSS 0.00446951f
c3 3 VSS 0.00456548f
c4 10 VSS 0.00204811f
c5 11 VSS 0.00209587f
c6 12 VSS 0.00209928f
c7 13 VSS 0.0198989f
r1 37 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r2 3 36 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r3 33 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3140 $Y=0.0675 $X2=0.3260 $Y2=0.0675
r4 12 33 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3140 $Y2=0.0675
r5 34 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 32 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r7 30 31 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r8 2 30 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.0675 $X2=0.2260 $Y2=0.0675
r9 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r10 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r11 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r12 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2180 $Y2=0.0360
r13 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r14 24 25 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2405
+ $Y=0.0360 $X2=0.2855 $Y2=0.0360
r15 23 24 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.0360 $X2=0.2405 $Y2=0.0360
r16 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.0360 $X2=0.2180 $Y2=0.0360
r17 21 22 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.0360 $X2=0.2090 $Y2=0.0360
r18 20 21 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1840
+ $Y=0.0360 $X2=0.1995 $Y2=0.0360
r19 19 20 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.0360 $X2=0.1840 $Y2=0.0360
r20 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1465 $Y2=0.0360
r21 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r22 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r23 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r24 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r25 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r26 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00532382f
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%NET22 VSS 15 18 31 34 37 38 12 2 3 11 10 1 13
c1 1 VSS 0.00452766f
c2 2 VSS 0.00459721f
c3 3 VSS 0.00433548f
c4 10 VSS 0.00209679f
c5 11 VSS 0.00208798f
c6 12 VSS 0.00204307f
c7 13 VSS 0.0190931f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0675 $X2=0.9865 $Y2=0.0675
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9720 $Y=0.0675 $X2=0.9865 $Y2=0.0675
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.0675 $X2=0.9720 $Y2=0.0675
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.0675 $X2=0.9575 $Y2=0.0675
r5 34 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r6 2 33 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.0675 $X2=0.8785 $Y2=0.0675
r7 30 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.0675 $X2=0.8660 $Y2=0.0675
r8 11 30 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.0675 $X2=0.8540 $Y2=0.0675
r9 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.0675 $X2=0.8495 $Y2=0.0675
r10 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9720 $Y=0.0675
+ $X2=0.9720 $Y2=0.0360
r11 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.0675
+ $X2=0.8605 $Y2=0.0360
r12 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9335
+ $Y=0.0360 $X2=0.9720 $Y2=0.0360
r13 26 27 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.9035
+ $Y=0.0360 $X2=0.9335 $Y2=0.0360
r14 25 26 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.0360 $X2=0.9035 $Y2=0.0360
r15 24 25 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8790
+ $Y=0.0360 $X2=0.8940 $Y2=0.0360
r16 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8695
+ $Y=0.0360 $X2=0.8790 $Y2=0.0360
r17 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8605
+ $Y=0.0360 $X2=0.8695 $Y2=0.0360
r18 21 22 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8395
+ $Y=0.0360 $X2=0.8605 $Y2=0.0360
r19 20 21 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7945
+ $Y=0.0360 $X2=0.8395 $Y2=0.0360
r20 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7945 $Y2=0.0360
r21 13 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.0360 $X2=0.7560 $Y2=0.0360
r22 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r23 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r24 16 17 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7660 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r25 1 16 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7540 $Y=0.0675 $X2=0.7660 $Y2=0.0675
r26 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7540 $Y2=0.0675
r27 15 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%B VSS 39 5 6 7 8 9 10 12 1 2 15 13 11 14
c1 1 VSS 0.0175768f
c2 2 VSS 0.0175017f
c3 5 VSS 0.0496508f
c4 6 VSS 0.0495767f
c5 7 VSS 0.0474882f
c6 8 VSS 0.0474156f
c7 9 VSS 0.0495767f
c8 10 VSS 0.0496424f
c9 11 VSS 0.00646803f
c10 12 VSS 0.0123004f
c11 13 VSS 0.00641336f
c12 14 VSS 0.00567405f
c13 15 VSS 0.0056573f
r1 5 52 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r2 6 46 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 7 56 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r4 54 56 2.38179 $w=2e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3485
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r5 50 52 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 49 50 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r7 47 49 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r8 46 47 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r9 44 46 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 43 44 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r11 41 54 3.87634 $w=1.88833e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3395 $Y=0.1350 $X2=0.3485 $Y2=0.1350
r12 1 41 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3370
+ $Y=0.1350 $X2=0.3395 $Y2=0.1350
r13 1 43 12.9528 $w=1.33e-08 $l=1.3e-08 $layer=LIG $thickness=4.8e-08 $X=0.3370
+ $Y=0.1350 $X2=0.3240 $Y2=0.1350
r14 39 40 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1350 $X2=0.3470 $Y2=0.1540
r15 39 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3470 $Y=0.1350
+ $X2=0.3485 $Y2=0.1350
r16 11 14 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3470 $Y=0.1765 $X2=0.3470 $Y2=0.1980
r17 11 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1765 $X2=0.3470 $Y2=0.1540
r18 14 37 22.7192 $w=1.34306e-08 $l=1.045e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.3470 $Y=0.1980 $X2=0.4515 $Y2=0.1980
r19 36 37 24.3683 $w=1.3e-08 $l=1.045e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.5560 $Y=0.1980 $X2=0.4515 $Y2=0.1980
r20 12 15 19.1048 $w=1.35056e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6450 $Y=0.1980 $X2=0.7340 $Y2=0.1980
r21 12 36 20.7539 $w=1.3e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6450
+ $Y=0.1980 $X2=0.5560 $Y2=0.1980
r22 15 35 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7340 $Y=0.1980 $X2=0.7340 $Y2=0.1765
r23 10 30 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r24 9 24 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r25 34 35 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.1540 $X2=0.7340 $Y2=0.1765
r26 33 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.1350 $X2=0.7340 $Y2=0.1540
r27 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.1170 $X2=0.7340 $Y2=0.1350
r28 13 32 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.1070 $X2=0.7340 $Y2=0.1170
r29 28 30 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8245 $Y=0.1350 $X2=0.8370 $Y2=0.1350
r30 27 28 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8100 $Y=0.1350 $X2=0.8245 $Y2=0.1350
r31 25 27 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7955 $Y=0.1350 $X2=0.8100 $Y2=0.1350
r32 24 25 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7955 $Y2=0.1350
r33 22 24 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1350 $X2=0.7830 $Y2=0.1350
r34 21 22 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1350 $X2=0.7705 $Y2=0.1350
r35 20 21 12.4546 $w=1.33e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7435 $Y=0.1350 $X2=0.7560 $Y2=0.1350
r36 19 20 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7410 $Y=0.1350 $X2=0.7435 $Y2=0.1350
r37 17 19 4.21574 $w=1.85111e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7320 $Y=0.1350 $X2=0.7410 $Y2=0.1350
r38 17 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7320 $Y=0.1350
+ $X2=0.7340 $Y2=0.1350
r39 2 17 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7220
+ $Y=0.1350 $X2=0.7320 $Y2=0.1350
r40 2 18 1.4509 $w=1.90429e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7220 $Y=0.1350 $X2=0.7185 $Y2=0.1350
r41 8 17 2.53767 $w=1.41765e-07 $l=3e-09 $layer=LIG $thickness=5.27059e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7320 $Y2=0.1350
r42 8 18 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7185 $Y2=0.1350
r43 8 19 2.3074 $w=1.91383e-07 $l=1.2e-08 $layer=LIG $thickness=5.46667e-08
+ $X=0.7290 $Y=0.1350 $X2=0.7410 $Y2=0.1350
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%C VSS 43 3 4 5 6 7 8 9 1
c1 1 VSS 0.0326239f
c2 3 VSS 0.0848729f
c3 4 VSS 0.0866439f
c4 5 VSS 0.0494061f
c5 6 VSS 0.0493875f
c6 7 VSS 0.0866524f
c7 8 VSS 0.0848742f
c8 9 VSS 0.00624413f
r1 8 41 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r2 3 35 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r3 4 29 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r4 5 23 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 43 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.1350 $X2=0.5560 $Y2=0.1160
r6 6 16 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r7 39 41 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r8 38 39 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r9 37 38 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r10 33 35 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r11 32 33 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r12 30 32 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r13 29 30 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r14 27 29 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r15 26 27 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r16 24 26 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r17 23 24 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r18 21 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r19 19 20 11.9564 $w=1.33e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5375 $Y=0.1350 $X2=0.5495 $Y2=0.1350
r20 19 21 11.9564 $w=1.33e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5375 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r21 17 20 4.98184 $w=1.33e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5545
+ $Y=0.1350 $X2=0.5495 $Y2=0.1350
r22 15 16 1.90543 $w=2e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.5710
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r23 14 15 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.5610
+ $Y=0.1350 $X2=0.5710 $Y2=0.1350
r24 14 17 3.76121 $w=1.74231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5610 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r25 43 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5560 $Y=0.1350
+ $X2=0.5610 $Y2=0.1350
r26 12 15 4.39635 $w=1.80294e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5795 $Y=0.1350 $X2=0.5710 $Y2=0.1350
r27 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5940 $Y=0.1350 $X2=0.5795 $Y2=0.1350
r28 10 11 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6085 $Y=0.1350 $X2=0.5940 $Y2=0.1350
r29 7 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r30 1 10 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6085 $Y2=0.1350
r31 1 37 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
r32 7 10 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6085 $Y2=0.1350
r33 7 37 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%A VSS 40 5 6 7 8 9 10 13 14 1 2 11 12 15
c1 1 VSS 0.00268717f
c2 2 VSS 0.00264513f
c3 5 VSS 0.00614987f
c4 6 VSS 0.00524015f
c5 7 VSS 0.0427219f
c6 8 VSS 0.0427119f
c7 9 VSS 0.00523818f
c8 10 VSS 0.00617432f
c9 11 VSS 0.00496212f
c10 12 VSS 0.00459602f
c11 13 VSS 0.00121296f
c12 14 VSS 0.00127972f
c13 15 VSS 0.095097f
r1 10 60 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r2 9 54 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1350
r3 8 47 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r4 58 60 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9865 $Y=0.1350 $X2=0.9990 $Y2=0.1350
r5 57 58 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9720 $Y=0.1350 $X2=0.9865 $Y2=0.1350
r6 55 57 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9575 $Y=0.1350 $X2=0.9720 $Y2=0.1350
r7 54 55 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9575 $Y2=0.1350
r8 52 54 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9325 $Y=0.1350 $X2=0.9450 $Y2=0.1350
r9 51 52 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9180 $Y=0.1350 $X2=0.9325 $Y2=0.1350
r10 50 51 13.451 $w=1.33e-08 $l=1.35e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9045 $Y=0.1350 $X2=0.9180 $Y2=0.1350
r11 49 50 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.9020 $Y=0.1350 $X2=0.9045 $Y2=0.1350
r12 46 47 2.54058 $w=2e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.8930
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r13 46 49 3.53695 $w=1.92556e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.8930 $Y=0.1350 $X2=0.9020 $Y2=0.1350
r14 2 46 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.8830
+ $Y=0.1350 $X2=0.8930 $Y2=0.1350
r15 14 44 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8940 $Y=0.1980 $X2=0.8940 $Y2=0.1845
r16 40 14 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8940 $Y=0.1890 $X2=0.8940
+ $Y2=0.1980
r17 43 44 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.1620 $X2=0.8940 $Y2=0.1845
r18 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.1350 $X2=0.8940 $Y2=0.1620
r19 42 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8940 $Y=0.1350
+ $X2=0.8930 $Y2=0.1350
r20 12 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.1170 $X2=0.8940 $Y2=0.1350
r21 40 44 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8940 $Y=0.1890 $X2=0.8940
+ $Y2=0.1845
r22 40 39 82.899 $w=1.3e-08 $l=3.555e-07 $layer=M2 $thickness=3.6e-08 $X=0.8940
+ $Y=0.1890 $X2=0.5385 $Y2=0.1890
r23 38 39 82.899 $w=1.3e-08 $l=3.555e-07 $layer=M2 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1890 $X2=0.5385 $Y2=0.1890
r24 15 38 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1715
+ $Y=0.1890 $X2=0.1830 $Y2=0.1890
r25 13 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1830 $Y=0.1980 $X2=0.1830 $Y2=0.1845
r26 13 38 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1830 $Y=0.1980 $X2=0.1830
+ $Y2=0.1890
r27 36 38 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1830 $Y=0.1845 $X2=0.1830
+ $Y2=0.1890
r28 35 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1620 $X2=0.1830 $Y2=0.1845
r29 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1350 $X2=0.1830 $Y2=0.1620
r30 11 34 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1160 $X2=0.1830 $Y2=0.1350
r31 7 31 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r32 6 23 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r33 29 31 2.06422 $w=2e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1855
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r34 29 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1855 $Y=0.1350
+ $X2=0.1830 $Y2=0.1350
r35 27 29 4.55514 $w=1.81389e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1855 $Y2=0.1350
r36 26 27 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r37 24 26 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r38 23 24 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r39 21 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r40 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r41 19 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r42 5 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r43 1 18 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r44 1 19 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r45 5 18 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r46 5 19 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_NAND3x2_ASAP7_75t_R%Y VSS 87 43 54 57 76 79 80 83 84 91 98 100 103 6
+ 2 3 7 35 25 28 1 8 27 33 37 29 32 36 34 26 31 4 5 30
c1 1 VSS 0.00413236f
c2 2 VSS 0.00292091f
c3 3 VSS 0.00765609f
c4 4 VSS 0.0100056f
c5 5 VSS 0.0097846f
c6 6 VSS 0.00291777f
c7 7 VSS 0.00777414f
c8 8 VSS 0.00412987f
c9 25 VSS 0.00234539f
c10 26 VSS 0.00217206f
c11 27 VSS 0.00217256f
c12 28 VSS 0.00233726f
c13 29 VSS 0.00347872f
c14 30 VSS 0.00472467f
c15 31 VSS 0.00471945f
c16 32 VSS 0.00346375f
c17 33 VSS 0.00283233f
c18 34 VSS 0.00211286f
c19 35 VSS 0.08904f
c20 36 VSS 0.00220201f
c21 37 VSS 0.00281372f
c22 38 VSS 0.00107557f
c23 39 VSS 0.00275985f
c24 40 VSS 0.00107557f
c25 41 VSS 0.00275985f
r1 103 102 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r2 101 102 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.0675 $X2=0.9325 $Y2=0.0675
r3 6 101 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.0675 $X2=0.9280 $Y2=0.0675
r4 27 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0675 $X2=0.9160 $Y2=0.0675
r5 100 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0675 $X2=0.9035 $Y2=0.0675
r6 28 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.0675 $X2=1.0240 $Y2=0.0675
r7 98 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.0675 $X2=1.0115 $Y2=0.0675
r8 6 95 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.0675
+ $X2=0.9180 $Y2=0.0720
r9 8 92 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.0675
+ $X2=1.0260 $Y2=0.0720
r10 95 96 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0720 $X2=0.9565 $Y2=0.0720
r11 92 93 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.0720 $X2=1.0395 $Y2=0.0720
r12 36 92 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.0015
+ $Y=0.0720 $X2=1.0260 $Y2=0.0720
r13 36 96 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0015
+ $Y=0.0720 $X2=0.9565 $Y2=0.0720
r14 40 89 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0720 $X2=1.0530 $Y2=0.0945
r15 40 93 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0720 $X2=1.0395 $Y2=0.0720
r16 32 7 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2025 $X2=0.9160 $Y2=0.2025
r17 91 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2025 $X2=0.9035 $Y2=0.2025
r18 87 88 5.42166 $w=1.3e-08 $l=2.32e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1430 $X2=1.0530 $Y2=0.1662
r19 87 86 4.13912 $w=1.3e-08 $l=1.78e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1430 $X2=1.0530 $Y2=0.1252
r20 86 89 7.17059 $w=1.3e-08 $l=3.07e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1252 $X2=1.0530 $Y2=0.0945
r21 85 88 7.40378 $w=1.3e-08 $l=3.18e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1980 $X2=1.0530 $Y2=0.1662
r22 37 41 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2160 $X2=1.0530 $Y2=0.2340
r23 37 85 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.2160 $X2=1.0530 $Y2=0.1980
r24 84 82 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r25 5 82 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r26 31 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2025 $X2=0.7020 $Y2=0.2025
r27 83 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2025 $X2=0.6875 $Y2=0.2025
r28 80 78 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r29 4 78 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r30 30 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r31 79 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r32 76 75 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r33 29 75 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r34 7 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2025
+ $X2=0.9180 $Y2=0.2340
r35 41 74 14.0912 $w=1.36667e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=0.9855 $Y2=0.2340
r36 5 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2025
+ $X2=0.7020 $Y2=0.2340
r37 4 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r38 3 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r39 73 74 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.2340 $X2=0.9855 $Y2=0.2340
r40 72 73 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9065
+ $Y=0.2340 $X2=0.9180 $Y2=0.2340
r41 71 72 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.9035
+ $Y=0.2340 $X2=0.9065 $Y2=0.2340
r42 70 71 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8845
+ $Y=0.2340 $X2=0.9035 $Y2=0.2340
r43 69 70 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8450
+ $Y=0.2340 $X2=0.8845 $Y2=0.2340
r44 68 69 14.3412 $w=1.3e-08 $l=6.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7835
+ $Y=0.2340 $X2=0.8450 $Y2=0.2340
r45 67 68 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7270
+ $Y=0.2340 $X2=0.7835 $Y2=0.2340
r46 66 67 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.2340 $X2=0.7270 $Y2=0.2340
r47 65 66 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.7020 $Y2=0.2340
r48 64 65 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r49 63 64 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r50 62 63 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3535 $Y2=0.2340
r51 61 62 14.8076 $w=1.3e-08 $l=6.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r52 60 61 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1925
+ $Y=0.2340 $X2=0.2335 $Y2=0.2340
r53 59 60 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1725
+ $Y=0.2340 $X2=0.1925 $Y2=0.2340
r54 58 59 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1725 $Y2=0.2340
r55 35 58 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r56 35 39 14.0912 $w=1.36667e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r57 39 52 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r58 57 56 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r59 2 56 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r60 53 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.0675 $X2=0.1640 $Y2=0.0675
r61 26 53 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1520 $Y2=0.0675
r62 54 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r63 51 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r64 50 51 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1475 $X2=0.0270 $Y2=0.1980
r65 33 38 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0935 $X2=0.0270 $Y2=0.0720
r66 33 50 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0935 $X2=0.0270 $Y2=0.1475
r67 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0720
r68 46 47 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.0720 $X2=0.1620 $Y2=0.0720
r69 45 46 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0785
+ $Y=0.0720 $X2=0.1235 $Y2=0.0720
r70 44 45 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0720 $X2=0.0785 $Y2=0.0720
r71 34 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0720 $X2=0.0540 $Y2=0.0720
r72 34 38 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0720 $X2=0.0270 $Y2=0.0720
r73 1 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0720
r74 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r75 25 42 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r76 3 29 1e-05
r77 1 25 1e-05
.ends


*
.SUBCKT NAND3x2_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0@4 N_MM0@4_d N_MM0@4_g N_MM0@4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@6 N_MM0@6_d N_MM0@6_g N_MM0@6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@5 N_MM0@5_d N_MM3_g N_MM0@5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@4 N_MM1@4_d N_MM1@4_g N_MM1@4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@6 N_MM1@6_d N_MM1@6_g N_MM1@6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@5 N_MM1@5_d N_MM4_g N_MM1@5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@6 N_MM2@6_d N_MM2@6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@5 N_MM2@5_d N_MM2@5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@4 N_MM2@4_d N_MM2@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@3 N_MM2@3_d N_MM2@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@3 N_MM1@3_d N_MM1@3_g N_MM1@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 N_MM0@3_d N_MM0@3_g N_MM0@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g N_MM0@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NAND3x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND3x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND3x2_ASAP7_75t_R%NET21 VSS N_MM2@3_d N_MM2@4_d N_MM2@6_d N_MM2@5_d
+ N_MM1@5_s N_MM2_d N_MM1@4_s N_MM1@6_s N_MM2@2_d N_MM1_s N_MM1@3_s N_MM1@2_s
+ N_NET21_24 N_NET21_20 N_NET21_4 N_NET21_19 N_NET21_5 N_NET21_2 N_NET21_1
+ N_NET21_6 N_NET21_25 N_NET21_23 N_NET21_22 N_NET21_3 N_NET21_21
+ PM_NAND3x2_ASAP7_75t_R%NET21
cc_1 N_NET21_24 N_B_1 0.000351528f
cc_2 N_NET21_24 N_B_2 0.00345866f
cc_3 N_NET21_24 N_MM1_g 0.000427521f
cc_4 N_NET21_20 N_MM4_g 0.0330829f
cc_5 N_NET21_4 N_B_12 0.000755578f
cc_6 N_NET21_19 N_MM1@4_g 0.0480323f
cc_7 N_NET21_5 N_MM1_g 0.00088448f
cc_8 N_NET21_2 N_MM4_g 0.000890729f
cc_9 N_NET21_1 N_MM1@4_g 0.00164785f
cc_10 N_NET21_6 N_MM1@3_g 0.00165125f
cc_11 N_NET21_19 N_B_1 0.00313053f
cc_12 N_NET21_25 N_B_13 0.00369785f
cc_13 N_NET21_25 N_B_11 0.00380495f
cc_14 N_NET21_23 N_MM1_g 0.0325408f
cc_15 N_NET21_24 N_MM1@2_g 0.0180669f
cc_16 N_NET21_19 N_MM1@6_g 0.018182f
cc_17 N_NET21_24 N_MM1@3_g 0.0489296f
cc_18 N_NET21_2 N_MM2@6_g 0.000673367f
cc_19 N_NET21_5 N_MM2@2_g 0.000683691f
cc_20 N_NET21_22 N_MM2@4_g 0.0482046f
cc_21 N_NET21_25 N_C_9 0.00165559f
cc_22 N_NET21_3 N_MM2@6_g 0.00168616f
cc_23 N_NET21_4 N_MM2@4_g 0.00173644f
cc_24 N_NET21_25 N_C_1 0.00241731f
cc_25 N_NET21_21 N_C_1 0.00635211f
cc_26 N_NET21_20 N_MM5_g 0.0325608f
cc_27 N_NET21_23 N_MM2@2_g 0.0326351f
cc_28 N_NET21_21 N_MM2@5_g 0.0181205f
cc_29 N_NET21_22 N_MM2@3_g 0.0181492f
cc_30 N_NET21_21 N_MM2@6_g 0.0498434f
cc_31 N_NET21_1 N_NET22__2_13 0.000719986f
cc_32 N_NET21_19 N_NET22__2_11 0.00110862f
cc_33 N_NET21_19 N_NET22__2_12 0.00110878f
cc_34 N_NET21_2 N_NET22__2_3 0.00122536f
cc_35 N_NET21_1 N_NET22__2_3 0.00309832f
cc_36 N_NET21_1 N_NET22__2_2 0.00418951f
cc_37 N_NET21_25 N_NET22__2_13 0.0111142f
x_PM_NAND3x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND3x2_ASAP7_75t_R%noxref_10
cc_38 N_noxref_10_1 N_MM0@4_g 0.00166515f
cc_39 N_noxref_10_1 N_Y_33 0.000257181f
cc_40 N_noxref_10_1 N_Y_1 0.000493806f
cc_41 N_noxref_10_1 N_Y_25 0.0366693f
x_PM_NAND3x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NAND3x2_ASAP7_75t_R%noxref_11
cc_42 N_noxref_11_1 N_MM0@4_g 0.00943298f
cc_43 N_noxref_11_1 N_Y_35 0.000119503f
cc_44 N_noxref_11_1 N_Y_33 0.000512236f
cc_45 N_noxref_11_1 N_Y_25 0.00154687f
cc_46 N_noxref_11_1 N_noxref_10_1 0.00194147f
x_PM_NAND3x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NAND3x2_ASAP7_75t_R%noxref_13
cc_47 N_noxref_13_1 N_MM0@2_g 0.00941492f
cc_48 N_noxref_13_1 N_Y_35 0.000120038f
cc_49 N_noxref_13_1 N_Y_37 0.000519266f
cc_50 N_noxref_13_1 N_Y_28 0.00156386f
cc_51 N_noxref_13_1 N_noxref_12_1 0.00193959f
x_PM_NAND3x2_ASAP7_75t_R%NET22__2 VSS N_MM0@4_s N_MM0@6_s N_MM0@5_s N_MM1@4_d
+ N_MM1@6_d N_MM1@5_d N_NET22__2_10 N_NET22__2_2 N_NET22__2_1 N_NET22__2_11
+ N_NET22__2_12 N_NET22__2_3 N_NET22__2_13 PM_NAND3x2_ASAP7_75t_R%NET22__2
cc_52 N_NET22__2_10 N_A_15 0.000298542f
cc_53 N_NET22__2_10 N_MM3_g 0.000450427f
cc_54 N_NET22__2_10 N_A_11 0.0010229f
cc_55 N_NET22__2_2 N_MM3_g 0.000999432f
cc_56 N_NET22__2_1 N_MM0@4_g 0.00165394f
cc_57 N_NET22__2_10 N_A_1 0.00268075f
cc_58 N_NET22__2_11 N_MM3_g 0.0327222f
cc_59 N_NET22__2_10 N_MM0@6_g 0.0181259f
cc_60 N_NET22__2_10 N_MM0@4_g 0.0484154f
cc_61 N_NET22__2_12 N_MM1@4_g 0.0011441f
cc_62 N_NET22__2_3 N_MM1@6_g 0.00183242f
cc_63 N_NET22__2_12 N_B_1 0.00280991f
cc_64 N_NET22__2_11 N_MM1@4_g 0.0326023f
cc_65 N_NET22__2_12 N_MM4_g 0.0180651f
cc_66 N_NET22__2_12 N_MM1@6_g 0.0487545f
x_PM_NAND3x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NAND3x2_ASAP7_75t_R%noxref_12
cc_67 N_noxref_12_1 N_MM0@2_g 0.00166475f
cc_68 N_noxref_12_1 N_Y_37 0.00026231f
cc_69 N_noxref_12_1 N_Y_8 0.000493689f
cc_70 N_noxref_12_1 N_Y_28 0.036689f
x_PM_NAND3x2_ASAP7_75t_R%NET22 VSS N_MM1_d N_MM1@3_d N_MM1@2_d N_MM0_s
+ N_MM0@3_s N_MM0@2_s N_NET22_12 N_NET22_2 N_NET22_3 N_NET22_11 N_NET22_10
+ N_NET22_1 N_NET22_13 PM_NAND3x2_ASAP7_75t_R%NET22
cc_71 N_NET22_12 N_A_15 0.000288357f
cc_72 N_NET22_12 N_MM0_g 0.000419353f
cc_73 N_NET22_12 N_A_12 0.000983601f
cc_74 N_NET22_2 N_MM0_g 0.00103575f
cc_75 N_NET22_3 N_MM0@3_g 0.00164114f
cc_76 N_NET22_12 N_A_2 0.00268213f
cc_77 N_NET22_11 N_MM0_g 0.0326717f
cc_78 N_NET22_12 N_MM0@2_g 0.0180858f
cc_79 N_NET22_12 N_MM0@3_g 0.0483812f
cc_80 N_NET22_10 N_MM1@2_g 0.00114222f
cc_81 N_NET22_1 N_MM1_g 0.00180501f
cc_82 N_NET22_10 N_B_2 0.00277151f
cc_83 N_NET22_11 N_MM1@2_g 0.0325529f
cc_84 N_NET22_10 N_MM1@3_g 0.0181542f
cc_85 N_NET22_10 N_MM1_g 0.0485581f
cc_86 N_NET22_13 N_NET21_6 0.000804942f
cc_87 N_NET22_10 N_NET21_24 0.00110937f
cc_88 N_NET22_10 N_NET21_23 0.00111001f
cc_89 N_NET22_2 N_NET21_6 0.00139686f
cc_90 N_NET22_1 N_NET21_6 0.00281538f
cc_91 N_NET22_1 N_NET21_5 0.00434741f
cc_92 N_NET22_13 N_NET21_25 0.01076f
x_PM_NAND3x2_ASAP7_75t_R%B VSS B N_MM1@4_g N_MM1@6_g N_MM4_g N_MM1_g N_MM1@3_g
+ N_MM1@2_g N_B_12 N_B_1 N_B_2 N_B_15 N_B_13 N_B_11 N_B_14
+ PM_NAND3x2_ASAP7_75t_R%B
cc_93 N_B_12 N_A_13 8.97689e-20
cc_94 N_B_12 N_A_14 9.52626e-20
cc_95 N_B_12 N_A_1 9.78146e-20
cc_96 N_B_12 N_A_2 0.000108273f
cc_97 N_B_1 N_A_11 0.000219391f
cc_98 N_B_2 N_A_12 0.000229061f
cc_99 N_B_15 N_A_15 0.000317199f
cc_100 N_B_13 N_A_15 0.00106103f
cc_101 N_B_11 N_A_15 0.0011086f
cc_102 N_B_2 N_A_2 0.00115345f
cc_103 N_B_1 N_A_1 0.00117698f
cc_104 N_MM1@2_g N_MM0_g 0.00341735f
cc_105 N_MM1@4_g N_MM3_g 0.00341994f
cc_106 N_B_14 N_A_15 0.00389114f
cc_107 N_B_12 N_A_15 0.00847259f
x_PM_NAND3x2_ASAP7_75t_R%C VSS C N_MM5_g N_MM2@6_g N_MM2@5_g N_MM2@4_g
+ N_MM2@3_g N_MM2@2_g N_C_9 N_C_1 PM_NAND3x2_ASAP7_75t_R%C
cc_108 N_C_9 N_B_13 0.000173318f
cc_109 N_C_9 N_B_1 0.000352602f
cc_110 N_C_9 N_B_2 0.000355509f
cc_111 N_C_1 N_B_12 0.00266199f
cc_112 N_MM2@2_g N_MM1_g 0.00340201f
cc_113 N_MM5_g N_MM4_g 0.00340573f
cc_114 N_C_9 N_B_12 0.00663854f
x_PM_NAND3x2_ASAP7_75t_R%A VSS A N_MM0@4_g N_MM0@6_g N_MM3_g N_MM0_g N_MM0@3_g
+ N_MM0@2_g N_A_13 N_A_14 N_A_1 N_A_2 N_A_11 N_A_12 N_A_15
+ PM_NAND3x2_ASAP7_75t_R%A
x_PM_NAND3x2_ASAP7_75t_R%Y VSS Y N_MM0@4_d N_MM0@6_d N_MM0@5_d N_MM3_d N_MM4_d
+ N_MM5_d N_MM5@2_d N_MM4@2_d N_MM3@2_d N_MM0@2_d N_MM0_d N_MM0@3_d N_Y_6 N_Y_2
+ N_Y_3 N_Y_7 N_Y_35 N_Y_25 N_Y_28 N_Y_1 N_Y_8 N_Y_27 N_Y_33 N_Y_37 N_Y_29
+ N_Y_32 N_Y_36 N_Y_34 N_Y_26 N_Y_31 N_Y_4 N_Y_5 N_Y_30 PM_NAND3x2_ASAP7_75t_R%Y
cc_115 N_Y_6 N_A_12 0.000252815f
cc_116 N_Y_2 N_A_11 0.000270527f
cc_117 N_Y_3 N_A_13 0.000331069f
cc_118 N_Y_7 N_A_14 0.000331232f
cc_119 N_Y_35 N_A_12 0.000344087f
cc_120 N_Y_35 N_A_11 0.000361641f
cc_121 N_Y_25 N_MM0@4_g 0.0353043f
cc_122 N_Y_28 N_MM0@2_g 0.0353211f
cc_123 N_Y_2 N_A_1 0.000596651f
cc_124 N_Y_6 N_A_2 0.000609278f
cc_125 N_Y_1 N_MM0@4_g 0.000838297f
cc_126 N_Y_8 N_MM0@2_g 0.000840601f
cc_127 N_Y_27 N_MM0_g 0.0681987f
cc_128 N_Y_33 N_A_1 0.00104373f
cc_129 N_Y_37 N_A_2 0.00107387f
cc_130 N_Y_29 N_MM3_g 0.0119451f
cc_131 N_Y_32 N_MM0_g 0.0330825f
cc_132 N_Y_36 N_A_2 0.00142223f
cc_133 N_Y_34 N_A_1 0.00152675f
cc_134 N_Y_7 N_A_12 0.00179944f
cc_135 N_Y_2 N_MM0@6_g 0.00188615f
cc_136 N_Y_6 N_MM0_g 0.00188692f
cc_137 N_Y_3 N_A_11 0.00202409f
cc_138 N_Y_35 N_A_14 0.002548f
cc_139 N_Y_35 N_A_13 0.00262913f
cc_140 N_Y_7 N_MM0_g 0.00288396f
cc_141 N_Y_3 N_MM0@6_g 0.00293367f
cc_142 N_Y_29 N_A_1 0.00633178f
cc_143 N_Y_32 N_A_2 0.00641257f
cc_144 N_Y_35 N_A_15 0.0171287f
cc_145 N_Y_29 N_MM0@6_g 0.0211879f
cc_146 N_Y_26 N_MM3_g 0.0372894f
cc_147 N_Y_27 N_MM0@3_g 0.0378379f
cc_148 N_Y_26 N_MM0@6_g 0.0691475f
cc_149 N_Y_31 N_MM4_g 0.00012362f
cc_150 N_Y_27 N_MM4_g 0.000146066f
cc_151 N_Y_26 N_MM4_g 0.000151843f
cc_152 N_Y_4 N_B_1 0.000184756f
cc_153 N_Y_5 N_B_2 0.00019088f
cc_154 N_Y_4 N_B_12 0.000426701f
cc_155 N_Y_31 N_MM1_g 0.0339905f
cc_156 N_Y_5 N_B_12 0.000449419f
cc_157 N_Y_5 N_B_13 0.000566814f
cc_158 N_Y_4 N_B_11 0.000597013f
cc_159 N_Y_30 N_B_1 0.00088808f
cc_160 N_Y_31 N_B_2 0.000957968f
cc_161 N_Y_4 N_MM4_g 0.00171126f
cc_162 N_Y_5 N_MM1_g 0.0017406f
cc_163 N_Y_35 N_B_15 0.00854168f
cc_164 N_Y_35 N_B_14 0.00877197f
cc_165 N_Y_35 N_B_12 0.0136897f
cc_166 N_Y_30 N_MM4_g 0.034475f
cc_167 N_Y_30 N_MM2@2_g 0.000590939f
cc_168 N_Y_35 N_MM2@2_g 0.000594092f
cc_169 N_Y_4 N_MM5_g 0.000696192f
cc_170 N_Y_5 N_MM2@2_g 0.000731564f
cc_171 N_Y_35 N_C_1 0.00149282f
cc_172 N_Y_30 N_MM5_g 0.0335408f
cc_173 N_Y_31 N_MM2@2_g 0.0345379f
cc_174 N_Y_33 N_NET22__2_13 0.000137094f
cc_175 N_Y_1 N_NET22__2_13 0.000202076f
cc_176 N_Y_2 N_NET22__2_13 0.000957144f
cc_177 N_Y_26 N_NET22__2_13 0.0005562f
cc_178 N_Y_25 N_NET22__2_13 0.000556796f
cc_179 N_Y_26 N_NET22__2_10 0.00110975f
cc_180 N_Y_25 N_NET22__2_10 0.00112075f
cc_181 N_Y_2 N_NET22__2_2 0.00133504f
cc_182 N_Y_2 N_NET22__2_1 0.00277702f
cc_183 N_Y_1 N_NET22__2_1 0.00454861f
cc_184 N_Y_34 N_NET22__2_13 0.00944555f
cc_185 N_Y_37 N_NET22_13 0.000128804f
cc_186 N_Y_6 N_NET22_13 0.000955501f
cc_187 N_Y_8 N_NET22_13 0.000261443f
cc_188 N_Y_28 N_NET22_13 0.000554196f
cc_189 N_Y_27 N_NET22_13 0.000554413f
cc_190 N_Y_27 N_NET22_11 0.00110908f
cc_191 N_Y_27 N_NET22_12 0.00111793f
cc_192 N_Y_8 N_NET22_3 0.00126235f
cc_193 N_Y_6 N_NET22_3 0.00327716f
cc_194 N_Y_6 N_NET22_2 0.00412757f
cc_195 N_Y_36 N_NET22_13 0.00942805f
*END of NAND3x2_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND3xp33_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND3xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND3xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND3xp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0328156f
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0425341f
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%NET21 VSS 2 3 1
c1 1 VSS 0.000895961f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%NET22 VSS 2 3 1
c1 1 VSS 0.000896488f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00496019f
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00377924f
c2 3 VSS 0.0715716f
c3 4 VSS 0.0161826f
r1 8 4 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0800
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0044853f
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%Y VSS 23 18 36 39 40 10 1 14 11 13 3 12
c1 1 VSS 0.00619571f
c2 3 VSS 0.00899941f
c3 10 VSS 0.00257521f
c4 11 VSS 0.0101278f
c5 12 VSS 0.00402507f
c6 13 VSS 0.00294191f
c7 14 VSS 0.0137099f
c8 15 VSS 0.00616722f
c9 16 VSS 0.00303517f
r1 40 38 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r2 3 38 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r3 12 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r4 39 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r5 36 35 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r6 11 35 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r7 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r8 11 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0000 $Y=0.0000
+ $X2=0.0540 $Y2=0.2340
r9 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r10 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r11 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r12 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r13 28 29 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r14 27 28 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0655
+ $Y=0.2340 $X2=0.0700 $Y2=0.2340
r15 26 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0655 $Y2=0.2340
r16 14 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r17 14 16 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r18 16 25 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r19 24 25 9.50248 $w=1.3e-08 $l=4.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1717 $X2=0.0270 $Y2=0.2125
r20 23 24 6.70421 $w=1.3e-08 $l=2.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1430 $X2=0.0270 $Y2=0.1717
r21 23 22 8.56972 $w=1.3e-08 $l=3.68e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1430 $X2=0.0270 $Y2=0.1062
r22 13 21 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r23 13 22 11.368 $w=1.3e-08 $l=4.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1062
r24 15 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r25 15 21 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r26 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r27 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r28 10 17 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r29 1 10 1e-05
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00400017f
c2 3 VSS 0.0353255f
c3 4 VSS 0.00697114f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NAND3xp33_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00546707f
c2 3 VSS 0.0347811f
c3 4 VSS 0.0045595f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends


*
.SUBCKT NAND3xp33_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 N_MM5_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND3xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND3xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND3xp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NAND3xp33_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM2_g 0.00376529f
cc_2 N_noxref_12_1 N_noxref_11_1 0.00192458f
x_PM_NAND3xp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NAND3xp33_ASAP7_75t_R%noxref_11
cc_3 N_noxref_11_1 N_MM2_g 0.00186147f
x_PM_NAND3xp33_ASAP7_75t_R%NET21 VSS N_MM1_s N_MM2_d N_NET21_1
+ PM_NAND3xp33_ASAP7_75t_R%NET21
cc_4 N_NET21_1 N_MM1_g 0.0173002f
cc_5 N_NET21_1 N_MM2_g 0.0172f
x_PM_NAND3xp33_ASAP7_75t_R%NET22 VSS N_MM0_s N_MM1_d N_NET22_1
+ PM_NAND3xp33_ASAP7_75t_R%NET22
cc_6 N_NET22_1 N_MM0_g 0.0172597f
cc_7 N_NET22_1 N_MM1_g 0.0172392f
x_PM_NAND3xp33_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NAND3xp33_ASAP7_75t_R%noxref_9
cc_8 N_noxref_9_1 N_MM0_g 0.00160407f
cc_9 N_noxref_9_1 N_Y_10 0.0379529f
x_PM_NAND3xp33_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 N_C_4
+ PM_NAND3xp33_ASAP7_75t_R%C
cc_10 N_C_1 N_B_1 0.00142736f
cc_11 N_C_4 N_B_4 0.00638022f
cc_12 N_MM2_g N_MM1_g 0.00852254f
x_PM_NAND3xp33_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NAND3xp33_ASAP7_75t_R%noxref_10
cc_13 N_noxref_10_1 N_MM0_g 0.00350897f
cc_14 N_noxref_10_1 N_Y_11 0.0287215f
cc_15 N_noxref_10_1 N_noxref_9_1 0.00190033f
x_PM_NAND3xp33_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM3_d N_MM4_d N_MM5_d N_Y_10 N_Y_1
+ N_Y_14 N_Y_11 N_Y_13 N_Y_3 N_Y_12 PM_NAND3xp33_ASAP7_75t_R%Y
cc_16 N_Y_10 N_A_4 0.000513256f
cc_17 N_Y_1 N_A_1 0.00074937f
cc_18 N_Y_14 N_A_4 0.0010787f
cc_19 N_Y_10 N_A_1 0.00141958f
cc_20 N_Y_1 N_MM0_g 0.00171194f
cc_21 N_Y_11 N_MM0_g 0.0107795f
cc_22 N_Y_13 N_A_4 0.00811843f
cc_23 N_Y_10 N_MM0_g 0.0505647f
cc_24 N_Y_3 N_MM1_g 0.000708241f
cc_25 N_Y_14 N_B_4 0.00110952f
cc_26 N_Y_1 N_B_4 0.00205469f
cc_27 N_Y_12 N_MM1_g 0.0269214f
cc_28 N_Y_12 N_C_4 0.000650692f
cc_29 N_Y_3 N_C_4 0.00118493f
cc_30 N_Y_12 N_MM2_g 0.0262868f
x_PM_NAND3xp33_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4
+ PM_NAND3xp33_ASAP7_75t_R%B
cc_31 N_B_1 N_A_1 0.00163885f
cc_32 N_B_4 N_A_4 0.00573238f
cc_33 N_MM1_g N_MM0_g 0.00837908f
x_PM_NAND3xp33_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4
+ PM_NAND3xp33_ASAP7_75t_R%A
*END of NAND3xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND4xp25_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND4xp25_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND4xp25_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND4xp25_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0425498f
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%PD1 VSS 2 3 1
c1 1 VSS 0.000893243f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0053252f
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00495703f
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00452296f
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00497888f
c2 3 VSS 0.0345562f
c3 4 VSS 0.00428534f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%PD3 VSS 2 3 1
c1 1 VSS 0.000904734f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%PD2 VSS 2 3 1
c1 1 VSS 0.000835994f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%Y VSS 27 22 46 49 50 52 1 17 14 2 15 3 19 4 13
+ 16 18
c1 1 VSS 0.00759758f
c2 2 VSS 0.00840002f
c3 3 VSS 0.00614163f
c4 4 VSS 0.00682006f
c5 13 VSS 0.0025809f
c6 14 VSS 0.00338652f
c7 15 VSS 0.00391251f
c8 16 VSS 0.00314542f
c9 17 VSS 0.0231441f
c10 18 VSS 0.00289704f
c11 19 VSS 0.0059632f
c12 20 VSS 0.00306165f
r1 52 51 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r2 14 51 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r3 50 48 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 2 48 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 15 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r6 49 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r7 16 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r8 46 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r9 1 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2340
r10 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r11 4 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r12 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r17 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 36 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r19 35 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r20 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r21 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r22 32 33 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r23 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r24 17 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r25 17 32 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2540 $Y2=0.2340
r26 20 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2970 $Y2=0.2125
r27 20 31 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2835 $Y2=0.2340
r28 28 29 9.1527 $w=1.3e-08 $l=3.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1732 $X2=0.2970 $Y2=0.2125
r29 27 28 6.35442 $w=1.3e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1460 $X2=0.2970 $Y2=0.1732
r30 27 26 8.91951 $w=1.3e-08 $l=3.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1460 $X2=0.2970 $Y2=0.1077
r31 18 25 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r32 18 26 11.7178 $w=1.3e-08 $l=5.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.1077
r33 24 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r34 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r35 19 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r36 3 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r37 13 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r38 22 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r39 1 14 1e-05
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%D VSS 10 3 1 4
c1 1 VSS 0.00366781f
c2 3 VSS 0.0714432f
c3 4 VSS 0.015069f
r1 10 4 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0800
r2 7 9 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1350 $X2=0.0915 $Y2=0.1350
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r4 10 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 1 8 2.51167 $w=1.2975e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0695 $Y2=0.1350
r7 3 6 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r8 3 8 2.63307 $w=1.98865e-07 $l=1.15e-08 $layer=LIG $thickness=5.49565e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0695 $Y2=0.1350
r9 3 9 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1350
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00384407f
c2 3 VSS 0.0350364f
c3 4 VSS 0.00699143f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_NAND4xp25_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00435304f
c2 3 VSS 0.0356632f
c3 4 VSS 0.00741479f
r1 8 4 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0800
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends


*
.SUBCKT NAND4xp25_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND4xp25_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND4xp25_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND4xp25_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NAND4xp25_ASAP7_75t_R%noxref_11
cc_1 N_noxref_11_1 N_MM5_g 0.00185757f
x_PM_NAND4xp25_ASAP7_75t_R%PD1 VSS N_MM4_d N_MM0_s N_PD1_1
+ PM_NAND4xp25_ASAP7_75t_R%PD1
cc_2 N_PD1_1 N_MM4_g 0.0173348f
cc_3 N_PD1_1 N_MM0_g 0.0173963f
x_PM_NAND4xp25_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NAND4xp25_ASAP7_75t_R%noxref_12
cc_4 N_noxref_12_1 N_MM5_g 0.00373598f
cc_5 N_noxref_12_1 N_Y_14 0.0274378f
cc_6 N_noxref_12_1 N_noxref_11_1 0.00192378f
x_PM_NAND4xp25_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NAND4xp25_ASAP7_75t_R%noxref_13
cc_7 N_noxref_13_1 N_MM0_g 0.00159972f
cc_8 N_noxref_13_1 N_Y_13 0.0379798f
x_PM_NAND4xp25_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NAND4xp25_ASAP7_75t_R%noxref_14
cc_9 N_noxref_14_1 N_MM0_g 0.00351366f
cc_10 N_noxref_14_1 N_Y_16 0.0286735f
cc_11 N_noxref_14_1 N_noxref_13_1 0.00189464f
x_PM_NAND4xp25_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4
+ PM_NAND4xp25_ASAP7_75t_R%A
cc_12 N_A_1 N_B_1 0.00151116f
cc_13 N_A_4 N_B_4 0.00548571f
cc_14 N_MM0_g N_MM4_g 0.00837153f
x_PM_NAND4xp25_ASAP7_75t_R%PD3 VSS N_MM5_d N_MM3_s N_PD3_1
+ PM_NAND4xp25_ASAP7_75t_R%PD3
cc_15 N_PD3_1 N_MM5_g 0.0172283f
cc_16 N_PD3_1 N_MM3_g 0.0173833f
x_PM_NAND4xp25_ASAP7_75t_R%PD2 VSS N_MM3_d N_MM4_s N_PD2_1
+ PM_NAND4xp25_ASAP7_75t_R%PD2
cc_17 N_PD2_1 N_MM3_g 0.0172913f
cc_18 N_PD2_1 N_MM4_g 0.0173602f
x_PM_NAND4xp25_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM1_d N_MM6_d N_MM2_d N_MM7_d
+ N_Y_1 N_Y_17 N_Y_14 N_Y_2 N_Y_15 N_Y_3 N_Y_19 N_Y_4 N_Y_13 N_Y_16 N_Y_18
+ PM_NAND4xp25_ASAP7_75t_R%Y
cc_19 N_Y_1 N_MM5_g 0.000860044f
cc_20 N_Y_17 N_D_4 0.00133608f
cc_21 N_Y_1 N_D_4 0.00192806f
cc_22 N_Y_14 N_MM5_g 0.0256844f
cc_23 N_Y_2 N_MM3_g 0.000716385f
cc_24 N_Y_17 N_C_4 0.00118795f
cc_25 N_Y_2 N_C_4 0.00175319f
cc_26 N_Y_15 N_MM3_g 0.0255747f
cc_27 N_Y_3 N_MM4_g 0.000355127f
cc_28 N_Y_2 N_MM4_g 0.0007062f
cc_29 N_Y_17 N_B_4 0.00116085f
cc_30 N_Y_3 N_B_4 0.00208561f
cc_31 N_Y_15 N_MM4_g 0.0265088f
cc_32 N_Y_19 N_A_4 0.000524237f
cc_33 N_Y_3 N_A_1 0.0007369f
cc_34 N_Y_4 N_MM0_g 0.000768842f
cc_35 N_Y_17 N_A_4 0.00111798f
cc_36 N_Y_13 N_A_1 0.00120671f
cc_37 N_Y_3 N_MM0_g 0.00169564f
cc_38 N_Y_16 N_MM0_g 0.0107835f
cc_39 N_Y_18 N_A_4 0.00808856f
cc_40 N_Y_13 N_MM0_g 0.0498602f
x_PM_NAND4xp25_ASAP7_75t_R%D VSS D N_MM5_g N_D_1 N_D_4
+ PM_NAND4xp25_ASAP7_75t_R%D
x_PM_NAND4xp25_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4
+ PM_NAND4xp25_ASAP7_75t_R%B
cc_41 N_B_1 N_C_1 0.00148896f
cc_42 N_B_4 N_C_4 0.00645733f
cc_43 N_MM4_g N_MM3_g 0.00869632f
x_PM_NAND4xp25_ASAP7_75t_R%C VSS C N_MM3_g N_C_1 N_C_4
+ PM_NAND4xp25_ASAP7_75t_R%C
cc_44 N_C_1 N_D_1 0.00150061f
cc_45 N_C_4 N_D_4 0.00661377f
cc_46 N_MM3_g N_MM5_g 0.00856971f
*END of NAND4xp25_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND4xp75_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND4xp75_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND4xp75_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND4xp75_ASAP7_75t_R%PD2 VSS 16 17 29 30 33 34 10 13 1 11 12 3 2
c1 1 VSS 0.00300448f
c2 2 VSS 0.00310542f
c3 3 VSS 0.0030171f
c4 10 VSS 0.00209341f
c5 11 VSS 0.00206826f
c6 12 VSS 0.00204395f
c7 13 VSS 0.00316388f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r2 3 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r4 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r5 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r6 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r8 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r9 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4850 $Y2=0.0720
r10 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0720
r11 24 25 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.0720 $X2=0.4850 $Y2=0.0720
r12 23 24 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3995
+ $Y=0.0720 $X2=0.4440 $Y2=0.0720
r13 22 23 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0720 $X2=0.3995 $Y2=0.0720
r14 21 22 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3545
+ $Y=0.0720 $X2=0.3780 $Y2=0.0720
r15 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3230
+ $Y=0.0720 $X2=0.3545 $Y2=0.0720
r16 19 20 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2925
+ $Y=0.0720 $X2=0.3230 $Y2=0.0720
r17 18 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0720 $X2=0.2925 $Y2=0.0720
r18 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0720 $X2=0.2700 $Y2=0.0720
r19 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0720
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r22 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r23 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0420295f
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0322822f
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%PD3 VSS 16 17 28 29 32 33 10 1 11 12 3 13 2
c1 1 VSS 0.010125f
c2 2 VSS 0.00732217f
c3 3 VSS 0.0045847f
c4 10 VSS 0.00454305f
c5 11 VSS 0.00329064f
c6 12 VSS 0.00213687f
c7 13 VSS 0.0227397f
r1 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r2 3 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r4 32 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r5 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r6 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r8 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r9 3 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r10 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r11 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r12 22 23 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2405
+ $Y=0.0360 $X2=0.2855 $Y2=0.0360
r13 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2405 $Y2=0.0360
r14 20 21 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r15 19 20 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r16 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r17 13 18 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0935
+ $Y=0.0360 $X2=0.0970 $Y2=0.0360
r18 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r21 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r22 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00571266f
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0316126f
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%D VSS 28 3 4 5 1 9 8 11
c1 1 VSS 0.00936164f
c2 3 VSS 0.0704347f
c3 4 VSS 0.0700172f
c4 5 VSS 0.0697732f
c5 6 VSS 0.011871f
c6 7 VSS 0.0121691f
c7 8 VSS 0.00508237f
c8 9 VSS 0.0102698f
c9 10 VSS 0.00322956f
c10 11 VSS 0.0103509f
r1 11 38 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r2 9 37 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 7 10 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1720 $X2=0.0270 $Y2=0.1350
r4 7 38 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.2125
r5 36 37 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0665 $X2=0.0270 $Y2=0.0540
r6 35 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0945 $X2=0.0270 $Y2=0.0665
r7 6 10 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1225 $X2=0.0270 $Y2=0.1350
r8 6 35 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1225 $X2=0.0270 $Y2=0.0945
r9 10 30 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0465 $Y2=0.1350
r10 5 26 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r11 4 20 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r12 28 8 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0645 $Y2=0.1350
r13 8 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0645
+ $Y=0.1350 $X2=0.0465 $Y2=0.1350
r14 24 26 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r15 23 24 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r16 21 23 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r17 20 21 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r18 18 20 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r19 17 18 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r20 16 17 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r21 14 16 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r22 13 14 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r23 28 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r24 1 13 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r25 1 15 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r26 3 13 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r27 3 15 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r28 3 16 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%A VSS 21 3 4 5 1 6
c1 1 VSS 0.0151478f
c2 3 VSS 0.0383038f
c3 4 VSS 0.0382972f
c4 5 VSS 0.038381f
c5 6 VSS 0.00817684f
r1 5 18 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r2 3 12 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 21 20 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1225
r4 6 20 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1125 $X2=0.6210 $Y2=0.1225
r5 16 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r6 15 16 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r7 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r8 10 12 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5795 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r9 9 10 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.5940
+ $Y=0.1350 $X2=0.5795 $Y2=0.1350
r10 8 9 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.6085
+ $Y=0.1350 $X2=0.5940 $Y2=0.1350
r11 4 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r12 21 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
r13 4 8 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6085 $Y2=0.1350
r14 4 14 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%PD1 VSS 16 17 29 30 33 34 10 1 13 11 3 12 2
c1 1 VSS 0.00470933f
c2 2 VSS 0.00418586f
c3 3 VSS 0.00449437f
c4 10 VSS 0.00216508f
c5 11 VSS 0.00208556f
c6 12 VSS 0.00214848f
c7 13 VSS 0.0217837f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r2 1 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r3 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r4 33 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r5 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r6 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r8 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r9 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r10 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r11 25 26 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4700 $Y2=0.0360
r12 23 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5015
+ $Y=0.0360 $X2=0.4700 $Y2=0.0360
r13 22 23 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5175
+ $Y=0.0360 $X2=0.5015 $Y2=0.0360
r14 21 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5175 $Y2=0.0360
r15 20 21 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5645
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r16 13 18 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6095
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r17 13 20 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6095
+ $Y=0.0360 $X2=0.5645 $Y2=0.0360
r18 3 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r20 3 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r21 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6480 $Y2=0.0675
r22 16 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%B VSS 27 3 4 5 8 7 1 6
c1 1 VSS 0.0133489f
c2 3 VSS 0.0374324f
c3 4 VSS 0.0373087f
c4 5 VSS 0.0372892f
c5 6 VSS 0.00704484f
c6 7 VSS 0.00556692f
c7 8 VSS 0.00598963f
r1 8 29 1.30447 $w=1.47857e-08 $l=1.49833e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5400 $Y=0.1035 $X2=0.5265 $Y2=0.1100
r2 7 29 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1100 $X2=0.5265 $Y2=0.1100
r3 27 6 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1225
r4 6 7 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1225 $X2=0.5130 $Y2=0.1100
r5 5 22 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r6 4 15 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r7 27 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r8 21 22 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r9 19 21 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5035 $Y2=0.1350
r10 18 19 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r11 16 18 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r12 15 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r13 13 15 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r14 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r15 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r16 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r17 1 10 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r18 1 11 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r19 3 10 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r20 3 11 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%C VSS 7 3 4 5 8 1 6 9
c1 1 VSS 0.0119426f
c2 3 VSS 0.0367221f
c3 4 VSS 0.0368116f
c4 5 VSS 0.0368495f
c5 6 VSS 0.00541996f
c6 7 VSS 0.00655861f
c7 8 VSS 0.00598706f
c8 9 VSS 0.00496928f
r1 8 28 4.53284 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.1100 $X2=0.2405 $Y2=0.1100
r2 6 9 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1100 $X2=0.2970 $Y2=0.1100
r3 6 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1100 $X2=0.2405 $Y2=0.1100
r4 9 25 1.26576 $w=2.0056e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1100 $X2=0.2970 $Y2=0.1225
r5 5 22 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 7 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r7 7 25 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1225
r8 4 16 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 20 22 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r10 19 20 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r11 17 19 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r12 16 17 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r13 14 16 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r14 13 14 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r15 12 13 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r16 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r17 1 11 4.63801 $w=1.7681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r18 1 12 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r19 3 11 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r20 3 12 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NAND4xp75_ASAP7_75t_R%Y VSS 50 40 41 54 78 79 82 83 86 87 90 91 94
+ 95 98 99 33 28 1 2 27 3 29 5 31 4 30 34 26 6 32 8 35 7 25
c1 1 VSS 0.00877792f
c2 2 VSS 0.00878629f
c3 3 VSS 0.00872467f
c4 4 VSS 0.00848492f
c5 5 VSS 0.00814833f
c6 6 VSS 0.00280623f
c7 7 VSS 0.00814187f
c8 8 VSS 0.00414199f
c9 25 VSS 0.00210274f
c10 26 VSS 0.0023092f
c11 27 VSS 0.00396951f
c12 28 VSS 0.00391209f
c13 29 VSS 0.00389583f
c14 30 VSS 0.00385314f
c15 31 VSS 0.0038487f
c16 32 VSS 0.00379725f
c17 33 VSS 0.0571307f
c18 34 VSS 0.00175756f
c19 35 VSS 0.00374923f
c20 36 VSS 0.00105777f
c21 37 VSS 0.00338947f
r1 99 97 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 1 97 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 27 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 98 27 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 95 93 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r6 2 93 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r7 28 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r8 94 28 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r9 91 89 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2160 $X2=0.4465 $Y2=0.2160
r10 4 89 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2160 $X2=0.4465 $Y2=0.2160
r11 30 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2160 $X2=0.4320 $Y2=0.2160
r12 90 30 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2160 $X2=0.4175 $Y2=0.2160
r13 87 85 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r14 3 85 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2160 $X2=0.3385 $Y2=0.2160
r15 29 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2160 $X2=0.3240 $Y2=0.2160
r16 86 29 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2160 $X2=0.3095 $Y2=0.2160
r17 83 81 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2160 $X2=0.5545 $Y2=0.2160
r18 5 81 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2160 $X2=0.5545 $Y2=0.2160
r19 31 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2160 $X2=0.5400 $Y2=0.2160
r20 82 31 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2160 $X2=0.5255 $Y2=0.2160
r21 79 77 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2160 $X2=0.6625 $Y2=0.2160
r22 7 77 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.2160 $X2=0.6625 $Y2=0.2160
r23 32 7 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2160 $X2=0.6480 $Y2=0.2160
r24 78 32 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2160 $X2=0.6335 $Y2=0.2160
r25 1 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1080 $Y2=0.2340
r26 2 71 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r27 4 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2160
+ $X2=0.4320 $Y2=0.2340
r28 3 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2160
+ $X2=0.3240 $Y2=0.2340
r29 5 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2160
+ $X2=0.5400 $Y2=0.2340
r30 7 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2160
+ $X2=0.6480 $Y2=0.2340
r31 73 74 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r32 71 74 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r33 70 71 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r34 69 70 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r35 67 68 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4700 $Y2=0.2340
r36 66 67 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r37 65 66 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r38 64 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r39 64 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r40 63 68 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5015
+ $Y=0.2340 $X2=0.4700 $Y2=0.2340
r41 62 63 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5015 $Y2=0.2340
r42 61 62 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.2340 $X2=0.5130 $Y2=0.2340
r43 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5265 $Y2=0.2340
r44 59 60 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5645
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r45 58 59 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5960
+ $Y=0.2340 $X2=0.5645 $Y2=0.2340
r46 57 58 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.2340 $X2=0.5960 $Y2=0.2340
r47 55 56 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.2340 $X2=0.6885 $Y2=0.2340
r48 33 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.2340 $X2=0.6480 $Y2=0.2340
r49 33 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.2340 $X2=0.6210 $Y2=0.2340
r50 37 52 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.7290 $Y2=0.2125
r51 37 56 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.2340 $X2=0.6885 $Y2=0.2340
r52 26 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7000 $Y2=0.0675
r53 54 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r54 51 52 9.1527 $w=1.3e-08 $l=3.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1732 $X2=0.7290 $Y2=0.2125
r55 50 51 6.35442 $w=1.3e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1460 $X2=0.7290 $Y2=0.1732
r56 50 49 4.72209 $w=1.3e-08 $l=2.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1460 $X2=0.7290 $Y2=0.1257
r57 35 36 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0935 $X2=0.7290 $Y2=0.0720
r58 35 49 7.52037 $w=1.3e-08 $l=3.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0935 $X2=0.7290 $Y2=0.1257
r59 8 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0675
+ $X2=0.7030 $Y2=0.0720
r60 36 48 1.38235 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0720 $X2=0.7160 $Y2=0.0720
r61 47 48 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.7030
+ $Y=0.0720 $X2=0.7160 $Y2=0.0720
r62 46 47 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6800
+ $Y=0.0720 $X2=0.7030 $Y2=0.0720
r63 45 46 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0720 $X2=0.6800 $Y2=0.0720
r64 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0720 $X2=0.6480 $Y2=0.0720
r65 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6075
+ $Y=0.0720 $X2=0.6210 $Y2=0.0720
r66 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0720 $X2=0.6075 $Y2=0.0720
r67 34 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.0720 $X2=0.5940 $Y2=0.0720
r68 6 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0720
r69 40 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r70 6 39 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r71 25 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r72 41 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
.ends


*
.SUBCKT NAND4xp75_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 N_MM5@3_d N_MM7@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM7@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM6_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@3 N_MM3@3_d N_MM6@3_g N_MM3@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM6@2_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM2_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM2@3_g N_MM4@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM2@2_g N_MM4@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 N_MM0@3_d N_MM0@3_g N_MM0@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g N_MM0@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7@3 N_MM7@3_d N_MM7@3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7@2 N_MM7@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6@3 N_MM6@3_d N_MM6@3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM6@2 N_MM6@2_d N_MM6@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2@3 N_MM2@3_d N_MM2@3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2@2 N_MM2@2_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@3 N_MM1@3_d N_MM0@3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 N_MM1@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND4xp75_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND4xp75_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND4xp75_ASAP7_75t_R%PD2 VSS N_MM3_d N_MM3@3_d N_MM3@2_d N_MM4_s
+ N_MM4@3_s N_MM4@2_s N_PD2_10 N_PD2_13 N_PD2_1 N_PD2_11 N_PD2_12 N_PD2_3
+ N_PD2_2 PM_NAND4xp75_ASAP7_75t_R%PD2
cc_1 N_PD2_10 N_C_8 0.000482528f
cc_2 N_PD2_10 N_MM6@2_g 0.000726621f
cc_3 N_PD2_13 N_C_6 0.00166533f
cc_4 N_PD2_1 N_MM6_g 0.00187358f
cc_5 N_PD2_10 N_C_1 0.00290981f
cc_6 N_PD2_13 N_C_9 0.00408088f
cc_7 N_PD2_11 N_MM6@2_g 0.0325037f
cc_8 N_PD2_10 N_MM6@3_g 0.0180009f
cc_9 N_PD2_10 N_MM6_g 0.0491213f
cc_10 N_PD2_12 N_MM2_g 0.000739646f
cc_11 N_PD2_12 N_B_7 0.000776842f
cc_12 N_PD2_13 N_B_1 0.00154718f
cc_13 N_PD2_3 N_MM2@3_g 0.00179724f
cc_14 N_PD2_12 N_B_1 0.00363577f
cc_15 N_PD2_11 N_MM2_g 0.03253f
cc_16 N_PD2_12 N_MM2@2_g 0.0179415f
cc_17 N_PD2_12 N_MM2@3_g 0.0497524f
cc_18 N_PD2_10 N_PD3_13 0.00110098f
cc_19 N_PD2_10 N_PD3_11 0.00110427f
cc_20 N_PD2_2 N_PD3_3 0.00126023f
cc_21 N_PD2_1 N_PD3_3 0.00301881f
cc_22 N_PD2_1 N_PD3_2 0.00399239f
cc_23 N_PD2_13 N_PD3_13 0.0116848f
x_PM_NAND4xp75_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NAND4xp75_ASAP7_75t_R%noxref_11
cc_24 N_noxref_11_1 N_MM5_g 0.00247244f
x_PM_NAND4xp75_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NAND4xp75_ASAP7_75t_R%noxref_12
cc_25 N_noxref_12_1 N_MM5_g 0.00448205f
cc_26 N_noxref_12_1 N_noxref_11_1 0.00189547f
x_PM_NAND4xp75_ASAP7_75t_R%PD3 VSS N_MM5_d N_MM5@3_d N_MM5@2_d N_MM3_s
+ N_MM3@3_s N_MM3@2_s N_PD3_10 N_PD3_1 N_PD3_11 N_PD3_12 N_PD3_3 N_PD3_13
+ N_PD3_2 PM_NAND4xp75_ASAP7_75t_R%PD3
cc_27 N_PD3_10 N_MM7@2_g 0.00208827f
cc_28 N_PD3_10 N_D_9 0.000460643f
cc_29 N_PD3_1 N_MM5_g 0.00195338f
cc_30 N_PD3_10 N_D_1 0.00286924f
cc_31 N_PD3_11 N_MM7@2_g 0.032838f
cc_32 N_PD3_10 N_MM7@3_g 0.0181764f
cc_33 N_PD3_10 N_MM5_g 0.0494149f
cc_34 N_PD3_12 N_MM6_g 0.0018368f
cc_35 N_PD3_3 N_MM6@3_g 0.00184699f
cc_36 N_PD3_12 N_C_1 0.00259091f
cc_37 N_PD3_13 N_C_8 0.00308091f
cc_38 N_PD3_11 N_MM6_g 0.0328664f
cc_39 N_PD3_12 N_MM6@2_g 0.0180979f
cc_40 N_PD3_12 N_MM6@3_g 0.0496101f
x_PM_NAND4xp75_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NAND4xp75_ASAP7_75t_R%noxref_13
cc_41 N_noxref_13_1 N_MM0@2_g 0.00160127f
cc_42 N_noxref_13_1 N_Y_8 0.000494622f
cc_43 N_noxref_13_1 N_Y_26 0.0366794f
x_PM_NAND4xp75_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NAND4xp75_ASAP7_75t_R%noxref_14
cc_44 N_noxref_14_1 N_MM0@2_g 0.00348273f
cc_45 N_noxref_14_1 N_Y_35 0.000356781f
cc_46 N_noxref_14_1 N_Y_32 0.00123437f
cc_47 N_noxref_14_1 N_noxref_13_1 0.00188936f
x_PM_NAND4xp75_ASAP7_75t_R%D VSS D N_MM5_g N_MM7@3_g N_MM7@2_g N_D_1 N_D_9
+ N_D_8 N_D_11 PM_NAND4xp75_ASAP7_75t_R%D
x_PM_NAND4xp75_ASAP7_75t_R%A VSS A N_MM1_g N_MM0@3_g N_MM0@2_g N_A_1 N_A_6
+ PM_NAND4xp75_ASAP7_75t_R%A
cc_48 N_A_1 N_B_8 0.00158986f
cc_49 N_MM1_g N_MM2@2_g 0.00753392f
x_PM_NAND4xp75_ASAP7_75t_R%PD1 VSS N_MM0@3_s N_MM0@2_s N_MM4@2_d N_MM0_s
+ N_MM4_d N_MM4@3_d N_PD1_10 N_PD1_1 N_PD1_13 N_PD1_11 N_PD1_3 N_PD1_12 N_PD1_2
+ PM_NAND4xp75_ASAP7_75t_R%PD1
cc_50 N_PD1_10 N_MM2@2_g 0.00141331f
cc_51 N_PD1_1 N_MM2_g 0.00172316f
cc_52 N_PD1_13 N_B_8 0.00249002f
cc_53 N_PD1_10 N_B_1 0.00304713f
cc_54 N_PD1_11 N_MM2@2_g 0.0329888f
cc_55 N_PD1_10 N_MM2@3_g 0.0182387f
cc_56 N_PD1_10 N_MM2_g 0.049942f
cc_57 N_PD1_3 N_MM0@3_g 0.00176231f
cc_58 N_PD1_12 N_A_1 0.00276463f
cc_59 N_PD1_11 N_MM1_g 0.0329711f
cc_60 N_PD1_12 N_MM0@2_g 0.0181928f
cc_61 N_PD1_12 N_MM0@3_g 0.0500594f
cc_62 N_PD1_10 N_PD2_11 0.00110362f
cc_63 N_PD1_10 N_PD2_12 0.00110475f
cc_64 N_PD1_2 N_PD2_3 0.00125866f
cc_65 N_PD1_1 N_PD2_3 0.00273379f
cc_66 N_PD1_1 N_PD2_2 0.00443381f
cc_67 N_PD1_13 N_PD2_13 0.0121875f
x_PM_NAND4xp75_ASAP7_75t_R%B VSS B N_MM2_g N_MM2@3_g N_MM2@2_g N_B_8 N_B_7
+ N_B_1 N_B_6 PM_NAND4xp75_ASAP7_75t_R%B
cc_68 N_MM2_g N_MM6@2_g 0.00711785f
x_PM_NAND4xp75_ASAP7_75t_R%C VSS C N_MM6_g N_MM6@3_g N_MM6@2_g N_C_8 N_C_1
+ N_C_6 N_C_9 PM_NAND4xp75_ASAP7_75t_R%C
cc_69 N_C_8 N_D_1 0.0014776f
cc_70 N_MM6_g N_MM7@2_g 0.00675473f
x_PM_NAND4xp75_ASAP7_75t_R%Y VSS Y N_MM0@3_d N_MM0_d N_MM0@2_d N_MM1@3_d
+ N_MM1@2_d N_MM2@2_d N_MM1_d N_MM6@3_d N_MM6@2_d N_MM2_d N_MM2@3_d N_MM7@2_d
+ N_MM6_d N_MM7_d N_MM7@3_d N_Y_33 N_Y_28 N_Y_1 N_Y_2 N_Y_27 N_Y_3 N_Y_29 N_Y_5
+ N_Y_31 N_Y_4 N_Y_30 N_Y_34 N_Y_26 N_Y_6 N_Y_32 N_Y_8 N_Y_35 N_Y_7 N_Y_25
+ PM_NAND4xp75_ASAP7_75t_R%Y
cc_71 N_Y_33 N_MM5_g 0.000334357f
cc_72 N_Y_28 N_MM5_g 0.000349766f
cc_73 N_Y_1 N_D_8 0.000380953f
cc_74 N_Y_33 N_D_11 0.000440369f
cc_75 N_Y_2 N_MM7@2_g 0.000524803f
cc_76 N_Y_33 N_MM7@2_g 0.00109042f
cc_77 N_Y_1 N_MM5_g 0.00117559f
cc_78 N_Y_27 N_D_1 0.00118293f
cc_79 N_Y_28 N_MM7@2_g 0.0240423f
cc_80 N_Y_27 N_MM7@3_g 0.0134138f
cc_81 N_Y_27 N_MM5_g 0.0360321f
cc_82 N_Y_3 N_MM6@3_g 0.00135594f
cc_83 N_Y_2 N_MM6@3_g 0.000491299f
cc_84 N_Y_28 N_MM6@3_g 0.000331724f
cc_85 N_Y_2 N_MM6_g 0.000591732f
cc_86 N_Y_29 N_C_1 0.0010748f
cc_87 N_Y_3 N_C 0.00213014f
cc_88 N_Y_33 N_C 0.00215922f
cc_89 N_Y_28 N_MM6_g 0.0239931f
cc_90 N_Y_29 N_MM6@2_g 0.0133896f
cc_91 N_Y_29 N_MM6@3_g 0.0359398f
cc_92 N_Y_5 N_MM2_g 0.000376001f
cc_93 N_Y_33 N_MM2_g 0.000182894f
cc_94 N_Y_31 N_MM2_g 0.000349771f
cc_95 N_Y_5 N_MM2@2_g 0.000755662f
cc_96 N_Y_4 N_MM2_g 0.00100924f
cc_97 N_Y_30 N_B_1 0.00125468f
cc_98 N_Y_34 N_B_8 0.00150003f
cc_99 N_Y_33 N_B_6 0.00179908f
cc_100 N_Y_5 N_B_6 0.00226643f
cc_101 N_Y_31 N_MM2@2_g 0.0241288f
cc_102 N_Y_30 N_MM2@3_g 0.0134369f
cc_103 N_Y_30 N_MM2_g 0.0359754f
cc_104 N_Y_31 N_MM1_g 0.0109218f
cc_105 N_Y_26 N_MM1_g 0.000471525f
cc_106 N_Y_6 N_MM1_g 0.00232747f
cc_107 N_Y_5 N_MM1_g 0.000530773f
cc_108 N_Y_32 N_MM0@3_g 0.022058f
cc_109 N_Y_8 N_MM0@2_g 0.000854843f
cc_110 N_Y_35 N_A_1 0.000903209f
cc_111 N_Y_7 N_MM0@3_g 0.00126461f
cc_112 N_Y_34 N_A_6 0.00163551f
cc_113 N_Y_33 N_A_6 0.00168467f
cc_114 N_Y_7 N_A_6 0.00401328f
cc_115 N_Y_25 N_A_1 0.00470226f
cc_116 N_Y_26 N_MM0@2_g 0.0471037f
cc_117 N_Y_25 N_MM0@3_g 0.0319114f
cc_118 N_Y_25 N_MM1_g 0.0633623f
cc_119 N_Y_6 N_PD1_13 0.000831692f
cc_120 N_Y_8 N_PD1_13 0.000242348f
cc_121 N_Y_26 N_PD1_13 0.00055549f
cc_122 N_Y_25 N_PD1_13 0.000567827f
cc_123 N_Y_25 N_PD1_11 0.00110975f
cc_124 N_Y_25 N_PD1_12 0.00112749f
cc_125 N_Y_8 N_PD1_3 0.00128985f
cc_126 N_Y_6 N_PD1_3 0.0031692f
cc_127 N_Y_6 N_PD1_2 0.00408638f
cc_128 N_Y_34 N_PD1_13 0.010105f
*END of NAND4xp75_ASAP7_75t_R.pxi
.ENDS
** Design:	NAND5xp2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NAND5xp2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NAND5xp2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NAND5xp2_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000867033f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%NET023 VSS 2 3 1
c1 1 VSS 0.000839305f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%NET024 VSS 2 3 1
c1 1 VSS 0.000876239f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0327638f
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0425156f
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.0008834f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%D VSS 8 3 1 4
c1 1 VSS 0.00434955f
c2 3 VSS 0.0356348f
c3 4 VSS 0.00766739f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1340 $X2=0.2430 $Y2=0.0795
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1345
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1340
+ $X2=0.2430 $Y2=0.1345
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00504182f
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00458703f
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%E VSS 8 3 1 4
c1 1 VSS 0.00384861f
c2 3 VSS 0.0716212f
c3 4 VSS 0.0153107f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1340 $X2=0.2970 $Y2=0.0795
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1345
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1340
+ $X2=0.2970 $Y2=0.1345
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00396732f
c2 3 VSS 0.0351967f
c3 4 VSS 0.00714752f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1340 $X2=0.1890 $Y2=0.0795
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1345
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1345
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%A VSS 11 3 1 4
c1 1 VSS 0.00577627f
c2 3 VSS 0.0350661f
c3 4 VSS 0.00472551f
r1 11 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0810 $Y2=0.0975
r2 7 10 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1340 $X2=0.0915 $Y2=0.1340
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0905 $Y2=0.1340
r4 11 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1340
+ $X2=0.0810 $Y2=0.1340
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1340 $X2=0.0810 $Y2=0.1340
r6 1 8 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1340 $X2=0.0685 $Y2=0.1340
r7 3 6 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1340
r8 3 8 4.17867 $w=1.8386e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1340
r9 3 10 1.08747 $w=2.16729e-07 $l=1.05475e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1340
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%B VSS 10 3 1 4
c1 1 VSS 0.00418274f
c2 3 VSS 0.0351662f
c3 4 VSS 0.00703199f
r1 10 9 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.0975
r2 4 9 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0575 $X2=0.1350 $Y2=0.0975
r3 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1345
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1345
.ends

.subckt PM_NAND5xp2_ASAP7_75t_R%Y VSS 27 23 48 51 52 55 56 18 1 2 19 13 14 17 3
+ 15 4 16
c1 1 VSS 0.00591897f
c2 2 VSS 0.00683081f
c3 3 VSS 0.00843573f
c4 4 VSS 0.00862657f
c5 13 VSS 0.00254229f
c6 14 VSS 0.00313327f
c7 15 VSS 0.00389069f
c8 16 VSS 0.00402449f
c9 17 VSS 0.00266488f
c10 18 VSS 0.00418073f
c11 19 VSS 0.0277807f
c12 20 VSS 0.00259265f
c13 21 VSS 0.00288614f
r1 56 54 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r2 4 54 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r3 16 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2700 $Y2=0.2160
r4 55 16 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r5 52 50 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r6 3 50 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r7 15 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r8 51 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r9 48 47 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r10 14 47 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r11 4 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r12 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r13 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2340
r14 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r15 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r16 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r17 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r18 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r19 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r20 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r21 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r22 34 35 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r23 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r24 32 33 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0710
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r25 31 32 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0665
+ $Y=0.2340 $X2=0.0710 $Y2=0.2340
r26 30 31 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0665 $Y2=0.2340
r27 19 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r28 19 21 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.2340 $X2=0.0180 $Y2=0.2340
r29 21 29 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.2340 $X2=0.0180 $Y2=0.2125
r30 28 29 11.1348 $w=1.3e-08 $l=4.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1647 $X2=0.0180 $Y2=0.2125
r31 27 28 8.33653 $w=1.3e-08 $l=3.57e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1290 $X2=0.0180 $Y2=0.1647
r32 27 26 6.9374 $w=1.3e-08 $l=2.98e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.1290 $X2=0.0180 $Y2=0.0992
r33 17 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0180 $Y=0.0575 $X2=0.0180 $Y2=0.0360
r34 17 26 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.0180
+ $Y=0.0575 $X2=0.0180 $Y2=0.0992
r35 18 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r36 18 20 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0360
+ $Y=0.0360 $X2=0.0180 $Y2=0.0360
r37 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r38 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r39 13 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r40 2 14 1e-05
r41 1 13 1e-05
.ends


*
.SUBCKT NAND5xp2_ASAP7_75t_R VSS VDD A B C D E Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* E E
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 N_MM8_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NAND5xp2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NAND5xp2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NAND5xp2_ASAP7_75t_R%NET30 VSS N_MM3_s N_MM5_d N_NET30_1
+ PM_NAND5xp2_ASAP7_75t_R%NET30
cc_1 N_NET30_1 N_MM3_g 0.017451f
cc_2 N_NET30_1 N_MM5_g 0.0175574f
x_PM_NAND5xp2_ASAP7_75t_R%NET023 VSS N_MM4_s N_MM3_d N_NET023_1
+ PM_NAND5xp2_ASAP7_75t_R%NET023
cc_3 N_NET023_1 N_MM4_g 0.0174656f
cc_4 N_NET023_1 N_MM3_g 0.0175703f
x_PM_NAND5xp2_ASAP7_75t_R%NET024 VSS N_MM0_s N_MM4_d N_NET024_1
+ PM_NAND5xp2_ASAP7_75t_R%NET024
cc_5 N_NET024_1 N_MM0_g 0.0172216f
cc_6 N_NET024_1 N_MM4_g 0.017299f
x_PM_NAND5xp2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_NAND5xp2_ASAP7_75t_R%noxref_16
cc_7 N_noxref_16_1 N_MM6_g 0.00373938f
cc_8 N_noxref_16_1 N_noxref_15_1 0.0019191f
x_PM_NAND5xp2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_NAND5xp2_ASAP7_75t_R%noxref_15
cc_9 N_noxref_15_1 N_MM6_g 0.00185394f
x_PM_NAND5xp2_ASAP7_75t_R%NET29 VSS N_MM5_s N_MM6_d N_NET29_1
+ PM_NAND5xp2_ASAP7_75t_R%NET29
cc_10 N_NET29_1 N_MM5_g 0.0172631f
cc_11 N_NET29_1 N_MM6_g 0.017249f
x_PM_NAND5xp2_ASAP7_75t_R%D VSS D N_MM5_g N_D_1 N_D_4 PM_NAND5xp2_ASAP7_75t_R%D
cc_12 N_D_1 N_C_1 0.00169564f
cc_13 N_D_4 N_C_4 0.00669318f
cc_14 N_MM5_g N_MM3_g 0.00867162f
x_PM_NAND5xp2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NAND5xp2_ASAP7_75t_R%noxref_13
cc_15 N_noxref_13_1 N_MM0_g 0.00166732f
cc_16 N_noxref_13_1 N_Y_13 0.0379163f
x_PM_NAND5xp2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NAND5xp2_ASAP7_75t_R%noxref_14
cc_17 N_noxref_14_1 N_MM0_g 0.00359705f
cc_18 N_noxref_14_1 N_Y_14 0.0286439f
cc_19 N_noxref_14_1 N_noxref_13_1 0.00188773f
x_PM_NAND5xp2_ASAP7_75t_R%E VSS E N_MM6_g N_E_1 N_E_4 PM_NAND5xp2_ASAP7_75t_R%E
cc_20 N_E_1 N_D_1 0.00164564f
cc_21 N_E_4 N_D_4 0.00689455f
cc_22 N_MM6_g N_MM5_g 0.00849873f
x_PM_NAND5xp2_ASAP7_75t_R%C VSS C N_MM3_g N_C_1 N_C_4 PM_NAND5xp2_ASAP7_75t_R%C
cc_23 N_C_1 N_B_1 0.00165568f
cc_24 N_C_4 N_B_4 0.00637494f
cc_25 N_MM3_g N_MM4_g 0.00873726f
x_PM_NAND5xp2_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_NAND5xp2_ASAP7_75t_R%A
x_PM_NAND5xp2_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4 PM_NAND5xp2_ASAP7_75t_R%B
cc_26 N_B_1 N_A_1 0.00154357f
cc_27 N_B_4 N_A_4 0.00549913f
cc_28 N_MM4_g N_MM0_g 0.00840499f
x_PM_NAND5xp2_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM10_d N_MM2_d N_MM7_d N_MM8_d
+ N_MM9_d N_Y_18 N_Y_1 N_Y_2 N_Y_19 N_Y_13 N_Y_14 N_Y_17 N_Y_3 N_Y_15 N_Y_4
+ N_Y_16 PM_NAND5xp2_ASAP7_75t_R%Y
cc_29 N_Y_18 N_A_4 0.000543086f
cc_30 N_Y_1 N_A_1 0.000622361f
cc_31 N_Y_2 N_MM0_g 0.000785414f
cc_32 N_Y_19 N_A_4 0.0011933f
cc_33 N_Y_13 N_A_1 0.0017685f
cc_34 N_Y_1 N_MM0_g 0.00198435f
cc_35 N_Y_14 N_MM0_g 0.0106837f
cc_36 N_Y_17 N_A_4 0.00712421f
cc_37 N_Y_13 N_MM0_g 0.0498175f
cc_38 N_Y_1 N_MM4_g 0.000346737f
cc_39 N_Y_3 N_MM4_g 0.000671219f
cc_40 N_Y_19 N_B_4 0.00122756f
cc_41 N_Y_1 N_B_4 0.00204833f
cc_42 N_Y_15 N_MM4_g 0.026307f
cc_43 N_Y_3 N_MM3_g 0.000668277f
cc_44 N_Y_19 N_C_4 0.00122387f
cc_45 N_Y_3 N_C_4 0.0016857f
cc_46 N_Y_15 N_MM3_g 0.0255095f
cc_47 N_Y_4 N_MM5_g 0.000654399f
cc_48 N_Y_19 N_D_4 0.00120541f
cc_49 N_Y_4 N_D_4 0.00163859f
cc_50 N_Y_16 N_MM5_g 0.0253691f
cc_51 N_Y_4 N_MM6_g 0.000719657f
cc_52 N_Y_19 N_E_4 0.00115203f
cc_53 N_Y_4 N_E_4 0.00156067f
cc_54 N_Y_16 N_MM6_g 0.0253446f
*END of NAND5xp2_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR2x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR2x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR2x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR2x1_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00570428f
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00464577f
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00547517f
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00470074f
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%NET16 VSS 15 30 31 33 1 2 13 10 11 3 12
c1 1 VSS 0.00794623f
c2 2 VSS 0.00690454f
c3 3 VSS 0.0053913f
c4 10 VSS 0.00341366f
c5 11 VSS 0.00333528f
c6 12 VSS 0.00222771f
c7 13 VSS 0.0225349f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r8 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r9 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 24 25 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1865
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r11 23 24 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1865 $Y2=0.2340
r12 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r13 21 22 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r14 20 21 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1005
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r15 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0890
+ $Y=0.2340 $X2=0.1005 $Y2=0.2340
r16 18 19 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0735
+ $Y=0.2340 $X2=0.0890 $Y2=0.2340
r17 17 18 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0735 $Y2=0.2340
r18 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r19 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0500 $Y2=0.2340
r21 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r22 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r23 1 10 1e-05
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%B VSS 19 3 4 6 9 10 1 7 8
c1 1 VSS 0.00681184f
c2 3 VSS 0.0450362f
c3 4 VSS 0.00765883f
c4 5 VSS 0.00338132f
c5 6 VSS 0.00328272f
c6 7 VSS 0.00365899f
c7 8 VSS 0.0036217f
c8 9 VSS 0.00388731f
c9 10 VSS 0.00261675f
r1 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1350
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1980
r3 5 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1350
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r5 10 21 7.6809 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1730 $Y2=0.1350
r6 4 17 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r7 19 7 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2045 $Y2=0.1350
r8 7 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.1350 $X2=0.1730 $Y2=0.1350
r9 15 17 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r10 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r11 19 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2160 $Y=0.1350
+ $X2=0.2160 $Y2=0.1350
r12 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r13 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r14 1 12 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r15 1 13 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r16 3 12 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r17 3 13 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%A VSS 24 3 4 1 10 7
c1 1 VSS 0.00685814f
c2 3 VSS 0.0431718f
c3 4 VSS 0.080395f
c4 5 VSS 0.00919991f
c5 6 VSS 0.00474635f
c6 7 VSS 0.00219668f
c7 8 VSS 0.00891822f
c8 9 VSS 0.00235893f
c9 10 VSS 0.00409796f
r1 8 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 6 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r3 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1980
r4 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r6 5 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r7 9 26 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r8 24 7 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0580 $Y2=0.1350
r9 7 26 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0580
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 3 18 0.314665 $w=2.27e-07 $l=5e-10 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1355
r11 17 18 1.4198 $w=2.3e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.0850
+ $Y=0.1355 $X2=0.0810 $Y2=0.1355
r12 16 17 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1355 $X2=0.0850 $Y2=0.1355
r13 24 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1355
r14 14 17 2.56587 $w=2.10294e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1355 $X2=0.0850 $Y2=0.1355
r15 13 14 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1355 $X2=0.0935 $Y2=0.1355
r16 12 13 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1355 $X2=0.1080 $Y2=0.1355
r17 4 1 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1355
r18 1 12 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1355 $X2=0.1225 $Y2=0.1355
r19 1 23 2.59554 $w=2.2681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1355 $X2=0.1455 $Y2=0.1355
r20 4 12 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1355
r21 4 23 0.54388 $w=2.16967e-07 $l=1.05119e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1350 $Y=0.1350 $X2=0.1455 $Y2=0.1355
.ends

.subckt PM_NOR2x1_ASAP7_75t_R%Y VSS 31 19 28 40 43 13 10 1 2 11 15 3 14 12
c1 1 VSS 0.00790424f
c2 2 VSS 0.00773286f
c3 3 VSS 0.00288886f
c4 10 VSS 0.00351508f
c5 11 VSS 0.00343396f
c6 12 VSS 0.00210415f
c7 13 VSS 0.017967f
c8 14 VSS 0.000760453f
c9 15 VSS 0.0025081f
c10 16 VSS 0.00294593f
c11 17 VSS 0.000761443f
r1 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 41 42 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 3 41 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r4 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r5 40 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r6 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r7 37 38 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2275 $Y2=0.1980
r8 35 38 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2570
+ $Y=0.1980 $X2=0.2275 $Y2=0.1980
r9 14 17 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2860 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r10 14 35 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1980 $X2=0.2570 $Y2=0.1980
r11 17 34 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1665
r12 33 34 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1665
r13 32 33 2.15701 $w=1.3e-08 $l=9.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1257 $X2=0.2970 $Y2=0.1350
r14 31 32 0.174892 $w=1.3e-08 $l=7e-10 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1250 $X2=0.2970 $Y2=0.1257
r15 31 30 5.18847 $w=1.3e-08 $l=2.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1250 $X2=0.2970 $Y2=0.1027
r16 29 30 7.17059 $w=1.3e-08 $l=3.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.1027
r17 15 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0360
r18 15 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0720
r19 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r20 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r21 16 26 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2590 $Y2=0.0360
r22 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r23 25 26 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2275
+ $Y=0.0360 $X2=0.2590 $Y2=0.0360
r24 24 25 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2275 $Y2=0.0360
r25 23 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r26 22 23 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r27 21 22 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r28 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.0360 $X2=0.1120 $Y2=0.0360
r29 13 20 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0360 $X2=0.1030 $Y2=0.0360
r30 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r31 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r32 10 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r33 1 10 1e-05
.ends


*
.SUBCKT NOR2x1_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 VDD N_MM2_g N_MM3@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR2x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR2x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR2x1_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1 PM_NOR2x1_ASAP7_75t_R%noxref_8
cc_1 N_noxref_8_1 N_MM3_g 0.00245708f
cc_2 N_noxref_8_1 N_NET16_10 0.0363233f
cc_3 N_noxref_8_1 N_noxref_7_1 0.00192313f
x_PM_NOR2x1_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_NOR2x1_ASAP7_75t_R%noxref_9
cc_4 N_noxref_9_1 N_MM4@2_g 0.00905942f
cc_5 N_noxref_9_1 N_NET16_12 0.000647253f
cc_6 N_noxref_9_1 N_Y_11 0.00196246f
x_PM_NOR2x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR2x1_ASAP7_75t_R%noxref_10
cc_7 N_noxref_10_1 N_MM4@2_g 0.00163959f
cc_8 N_noxref_10_1 N_NET16_12 0.0364542f
cc_9 N_noxref_10_1 N_Y_12 0.000811132f
cc_10 N_noxref_10_1 N_noxref_9_1 0.00193647f
x_PM_NOR2x1_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1 PM_NOR2x1_ASAP7_75t_R%noxref_7
cc_11 N_noxref_7_1 N_MM3_g 0.0104974f
cc_12 N_noxref_7_1 N_NET16_10 0.00058955f
cc_13 N_noxref_7_1 N_Y_10 0.0005896f
x_PM_NOR2x1_ASAP7_75t_R%NET16 VSS N_MM3_s N_MM3@2_s N_MM4_d N_MM4@2_d N_NET16_1
+ N_NET16_2 N_NET16_13 N_NET16_10 N_NET16_11 N_NET16_3 N_NET16_12
+ PM_NOR2x1_ASAP7_75t_R%NET16
cc_14 N_NET16_1 N_MM3_g 0.00278629f
cc_15 N_NET16_2 N_MM2_g 0.000756787f
cc_16 N_NET16_13 N_MM2_g 0.00150598f
cc_17 N_NET16_13 N_A_10 0.00197364f
cc_18 N_NET16_10 N_A_1 0.0020573f
cc_19 N_NET16_11 N_MM2_g 0.0333652f
cc_20 N_NET16_10 N_MM3_g 0.0360029f
cc_21 N_NET16_2 N_MM4@2_g 0.000571509f
cc_22 N_NET16_3 N_MM4@2_g 0.000960428f
cc_23 N_NET16_2 N_MM1_g 0.00145907f
cc_24 N_NET16_12 N_B_1 0.00162816f
cc_25 N_NET16_13 N_B_9 0.00515139f
cc_26 N_NET16_11 N_MM1_g 0.0334917f
cc_27 N_NET16_12 N_MM4@2_g 0.0359084f
x_PM_NOR2x1_ASAP7_75t_R%B VSS B N_MM1_g N_MM4@2_g N_B_6 N_B_9 N_B_10 N_B_1
+ N_B_7 N_B_8 PM_NOR2x1_ASAP7_75t_R%B
cc_28 N_B_6 N_A_1 0.00061747f
cc_29 N_B_9 N_A_10 0.000634654f
cc_30 N_B_10 N_A_7 0.000992216f
cc_31 N_B_10 N_A_1 0.00163642f
cc_32 N_MM1_g N_MM2_g 0.00631947f
x_PM_NOR2x1_ASAP7_75t_R%A VSS A N_MM3_g N_MM2_g N_A_1 N_A_10 N_A_7
+ PM_NOR2x1_ASAP7_75t_R%A
x_PM_NOR2x1_ASAP7_75t_R%Y VSS Y N_MM2_s N_MM1_s N_MM4_s N_MM4@2_s N_Y_13 N_Y_10
+ N_Y_1 N_Y_2 N_Y_11 N_Y_15 N_Y_3 N_Y_14 N_Y_12 PM_NOR2x1_ASAP7_75t_R%Y
cc_33 N_Y_13 N_MM2_g 0.000543716f
cc_34 N_Y_10 N_A_1 0.00241857f
cc_35 N_Y_1 N_MM2_g 0.0024976f
cc_36 N_Y_10 N_MM3_g 0.0191439f
cc_37 N_Y_10 N_MM2_g 0.0537072f
cc_38 N_Y_1 N_MM4@2_g 0.000734626f
cc_39 N_Y_2 N_B_1 0.00100339f
cc_40 N_Y_11 N_MM1_g 0.0494042f
cc_41 N_Y_15 N_B_7 0.00120879f
cc_42 N_Y_3 N_MM4@2_g 0.00197408f
cc_43 N_Y_2 N_MM4@2_g 0.00252701f
cc_44 N_Y_14 N_B_7 0.00329365f
cc_45 N_Y_12 N_B_1 0.0048254f
cc_46 N_Y_13 N_B_8 0.00554488f
cc_47 N_Y_11 N_MM4@2_g 0.0212126f
cc_48 N_Y_12 N_MM4@2_g 0.0711161f
cc_49 N_Y_14 N_NET16_3 0.000685052f
cc_50 N_Y_12 N_NET16_12 0.0018404f
cc_51 N_Y_3 N_NET16_13 0.000790377f
cc_52 N_Y_15 N_NET16_3 0.00082016f
cc_53 N_Y_3 N_NET16_2 0.00139607f
cc_54 N_Y_3 N_NET16_3 0.00534593f
cc_55 N_Y_14 N_NET16_13 0.00988047f
*END of NOR2x1_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR2x1p5_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR2x1p5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR2x1p5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR2x1p5_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0419579f
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00517324f
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00523171f
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00467198f
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%A VSS 30 3 4 5 1 8
c1 1 VSS 0.012782f
c2 3 VSS 0.043499f
c3 4 VSS 0.0799274f
c4 5 VSS 0.0803303f
c5 6 VSS 0.0111119f
c6 7 VSS 0.0120162f
c7 8 VSS 0.00342554f
c8 9 VSS 0.00965413f
c9 10 VSS 0.00313796f
c10 11 VSS 0.0100487f
r1 11 37 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 9 35 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 7 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r5 7 36 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r6 34 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 6 34 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 10 32 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 5 28 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1355
r11 30 8 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0580 $Y2=0.1350
r12 8 32 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0580
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r13 3 19 0.314665 $w=2.27e-07 $l=5e-10 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1355
r14 26 28 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1355 $X2=0.1890 $Y2=0.1355
r15 25 26 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1355 $X2=0.1765 $Y2=0.1355
r16 24 25 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1355 $X2=0.1620 $Y2=0.1355
r17 18 19 1.4198 $w=2.3e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.0850
+ $Y=0.1355 $X2=0.0810 $Y2=0.1355
r18 17 18 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1355 $X2=0.0850 $Y2=0.1355
r19 30 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1355
r20 15 18 2.56587 $w=2.10294e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1355 $X2=0.0850 $Y2=0.1355
r21 14 15 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1355 $X2=0.0935 $Y2=0.1355
r22 13 14 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1355 $X2=0.1080 $Y2=0.1355
r23 4 1 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1355
r24 1 13 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1355 $X2=0.1225 $Y2=0.1355
r25 1 24 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1355 $X2=0.1475 $Y2=0.1355
r26 4 13 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1355
r27 4 24 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1355
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%NET16 VSS 17 20 35 36 38 41 11 1 12 13 2 3 15 14
c1 1 VSS 0.00935518f
c2 2 VSS 0.00749257f
c3 3 VSS 0.00284821f
c4 11 VSS 0.00439213f
c5 12 VSS 0.00319088f
c6 13 VSS 0.00207691f
c7 14 VSS 0.0121507f
c8 15 VSS 0.00155201f
r1 41 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 39 40 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 3 39 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.2025 $X2=0.3340 $Y2=0.2025
r4 13 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r5 38 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r6 3 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r7 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r8 2 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r9 12 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r10 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r11 30 31 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2880
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r12 29 30 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2590
+ $Y=0.1980 $X2=0.2880 $Y2=0.1980
r13 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2410
+ $Y=0.1980 $X2=0.2590 $Y2=0.1980
r14 27 28 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2410 $Y2=0.1980
r15 15 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r16 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r17 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r18 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r19 24 25 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1730
+ $Y=0.2340 $X2=0.2045 $Y2=0.2340
r20 23 24 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.2340 $X2=0.1730 $Y2=0.2340
r21 22 23 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r22 21 22 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.2340 $X2=0.1120 $Y2=0.2340
r23 14 21 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.2340 $X2=0.1030 $Y2=0.2340
r24 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1120 $Y2=0.2340
r25 20 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r26 1 19 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r27 16 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.2025 $X2=0.1100 $Y2=0.2025
r28 11 16 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.0980 $Y2=0.2025
r29 17 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%B VSS 33 3 4 5 7 6 8 11 9 1 10
c1 1 VSS 0.0124455f
c2 3 VSS 0.0460457f
c3 4 VSS 0.045594f
c4 5 VSS 0.00865404f
c5 6 VSS 0.00428271f
c6 7 VSS 0.00434276f
c7 8 VSS 0.00542429f
c8 9 VSS 0.00467486f
c9 10 VSS 0.00487546f
c10 11 VSS 0.00356222f
r1 7 34 5.62944 $w=1.37143e-08 $l=2.63e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1402
r2 7 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1665 $X2=0.1350 $Y2=0.1980
r3 6 11 5.73148 $w=1.38716e-08 $l=2.72e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1307
r4 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r5 33 34 0.433689 $w=1.8e-08 $l=4.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.1402
r6 33 11 0.535733 $w=1.8e-08 $l=5.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.1307
r7 5 26 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r8 4 20 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 33 31 2.26632 $w=7.16216e-09 $l=1.8527e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1360 $X2=0.1535 $Y2=0.1350
r10 30 31 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1825
+ $Y=0.1350 $X2=0.1535 $Y2=0.1350
r11 8 28 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r12 8 30 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1350 $X2=0.1825 $Y2=0.1350
r13 24 26 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r14 23 24 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r15 21 23 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r16 20 21 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r17 18 20 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r18 17 18 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r19 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r20 14 16 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2525 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r21 13 14 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2525 $Y2=0.1350
r22 13 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r23 1 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r24 1 15 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2325 $Y2=0.1350
r25 3 13 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r26 3 15 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r27 3 16 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NOR2x1p5_ASAP7_75t_R%Y VSS 49 27 41 42 44 58 60 63 2 21 1 16 17 3 20
+ 23 19 5 4 18 22
c1 1 VSS 0.00805615f
c2 2 VSS 0.0089917f
c3 3 VSS 0.00452572f
c4 4 VSS 0.00777672f
c5 5 VSS 0.00513622f
c6 16 VSS 0.00349093f
c7 17 VSS 0.00416572f
c8 18 VSS 0.00348198f
c9 19 VSS 0.00219505f
c10 20 VSS 0.00232842f
c11 21 VSS 0.0289618f
c12 22 VSS 0.0113416f
c13 23 VSS 0.00341902f
c14 24 VSS 0.00302963f
c15 25 VSS 0.0028402f
r1 63 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 3 62 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 59 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2600 $Y=0.2025 $X2=0.2720 $Y2=0.2025
r4 19 59 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2600 $Y2=0.2025
r5 60 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r6 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r7 58 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r8 3 55 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r9 5 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r10 55 56 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r11 53 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r12 22 53 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r13 22 56 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r14 25 52 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4050 $Y2=0.2160
r15 25 54 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.3915 $Y2=0.2340
r16 51 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1980 $X2=0.4050 $Y2=0.2160
r17 50 51 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1672 $X2=0.4050 $Y2=0.1980
r18 49 50 5.18847 $w=1.3e-08 $l=2.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1450 $X2=0.4050 $Y2=0.1672
r19 49 48 0.174892 $w=1.3e-08 $l=8e-10 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1450 $X2=0.4050 $Y2=0.1442
r20 47 48 2.15701 $w=1.3e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1442
r21 46 47 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1035 $X2=0.4050 $Y2=0.1350
r22 45 46 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0720 $X2=0.4050 $Y2=0.1035
r23 23 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0360
r24 23 45 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0720
r25 18 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r26 44 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r27 42 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r28 2 40 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r29 17 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r30 41 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r31 24 38 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3670 $Y2=0.0360
r32 4 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r33 2 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r34 37 38 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3355
+ $Y=0.0360 $X2=0.3670 $Y2=0.0360
r35 36 37 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3355 $Y2=0.0360
r36 35 36 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r37 34 35 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2410
+ $Y=0.0360 $X2=0.2860 $Y2=0.0360
r38 33 34 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2410 $Y2=0.0360
r39 32 33 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1850
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r40 31 32 9.44418 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1445
+ $Y=0.0360 $X2=0.1850 $Y2=0.0360
r41 30 31 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1445 $Y2=0.0360
r42 29 30 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r43 28 29 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.0360 $X2=0.1120 $Y2=0.0360
r44 21 28 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0360 $X2=0.1030 $Y2=0.0360
r45 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r46 27 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r47 16 26 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r48 1 16 1e-05
.ends


*
.SUBCKT NOR2x1p5_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 VSS N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 VSS N_MM1@2_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@3 VDD N_MM2_g N_MM3@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 VDD N_MM2@2_g N_MM3@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM1@2_g N_MM4@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR2x1p5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR2x1p5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR2x1p5_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NOR2x1p5_ASAP7_75t_R%noxref_8
cc_1 N_noxref_8_1 N_MM3_g 0.00257755f
cc_2 N_noxref_8_1 N_noxref_7_1 0.00192522f
x_PM_NOR2x1p5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR2x1p5_ASAP7_75t_R%noxref_10
cc_3 N_noxref_10_1 N_MM4@2_g 0.00163201f
cc_4 N_noxref_10_1 N_Y_20 0.0376193f
cc_5 N_noxref_10_1 N_noxref_9_1 0.00193531f
x_PM_NOR2x1p5_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NOR2x1p5_ASAP7_75t_R%noxref_7
cc_6 N_noxref_7_1 N_MM3_g 0.0105631f
cc_7 N_noxref_7_1 N_Y_16 0.000598204f
x_PM_NOR2x1p5_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NOR2x1p5_ASAP7_75t_R%noxref_9
cc_8 N_noxref_9_1 N_MM4@2_g 0.00903111f
cc_9 N_noxref_9_1 N_Y_18 0.00262207f
x_PM_NOR2x1p5_ASAP7_75t_R%A VSS A N_MM3_g N_MM2_g N_MM2@2_g N_A_1 N_A_8
+ PM_NOR2x1p5_ASAP7_75t_R%A
x_PM_NOR2x1p5_ASAP7_75t_R%NET16 VSS N_MM3_s N_MM3@3_s N_MM3@2_s N_MM4_d
+ N_MM4@3_d N_MM4@2_d N_NET16_11 N_NET16_1 N_NET16_12 N_NET16_13 N_NET16_2
+ N_NET16_3 N_NET16_15 N_NET16_14 PM_NOR2x1p5_ASAP7_75t_R%NET16
cc_10 N_NET16_11 N_MM2@2_g 0.000736019f
cc_11 N_NET16_1 N_MM2_g 0.00202011f
cc_12 N_NET16_11 N_A_1 0.00311469f
cc_13 N_NET16_12 N_MM2@2_g 0.0328379f
cc_14 N_NET16_11 N_MM3_g 0.0180992f
cc_15 N_NET16_11 N_MM2_g 0.0502422f
cc_16 N_NET16_13 N_B_9 0.000672185f
cc_17 N_NET16_2 N_MM1_g 0.0010234f
cc_18 N_NET16_3 N_MM4@2_g 0.00168074f
cc_19 N_NET16_13 N_B_1 0.00316599f
cc_20 N_NET16_15 N_B_8 0.00345929f
cc_21 N_NET16_14 N_B_9 0.00492036f
cc_22 N_NET16_12 N_MM1_g 0.0328844f
cc_23 N_NET16_13 N_MM1@2_g 0.0180834f
cc_24 N_NET16_13 N_MM4@2_g 0.0506617f
x_PM_NOR2x1p5_ASAP7_75t_R%B VSS B N_MM1_g N_MM1@2_g N_MM4@2_g N_B_7 N_B_6 N_B_8
+ N_B_11 N_B_9 N_B_1 N_B_10 PM_NOR2x1p5_ASAP7_75t_R%B
cc_25 N_B_7 N_A_1 0.000691326f
cc_26 N_B_6 N_A_1 0.000736676f
cc_27 N_B_8 N_A_1 0.000966369f
cc_28 N_B_11 N_A_8 0.00106665f
cc_29 N_B_11 N_A_1 0.00257453f
cc_30 N_MM1_g N_MM2@2_g 0.00794653f
x_PM_NOR2x1p5_ASAP7_75t_R%Y VSS Y N_MM2_s N_MM2@2_s N_MM1_s N_MM1@2_s N_MM4@2_s
+ N_MM4_s N_MM4@3_s N_Y_2 N_Y_21 N_Y_1 N_Y_16 N_Y_17 N_Y_3 N_Y_20 N_Y_23 N_Y_19
+ N_Y_5 N_Y_4 N_Y_18 N_Y_22 PM_NOR2x1p5_ASAP7_75t_R%Y
cc_31 N_Y_2 N_MM2_g 0.00035512f
cc_32 N_Y_21 N_MM2_g 0.000941104f
cc_33 N_Y_21 N_MM2@2_g 0.000653348f
cc_34 N_Y_1 N_MM2_g 0.00248246f
cc_35 N_Y_16 N_A_1 0.00252345f
cc_36 N_Y_17 N_MM2@2_g 0.0242651f
cc_37 N_Y_16 N_MM3_g 0.0191226f
cc_38 N_Y_16 N_MM2_g 0.0532162f
cc_39 N_Y_3 N_MM1@2_g 0.00234856f
cc_40 N_Y_20 N_MM1@2_g 0.000452438f
cc_41 N_Y_1 N_MM1@2_g 0.000603766f
cc_42 N_Y_1 N_B_10 0.000604346f
cc_43 N_Y_2 N_MM1_g 0.000643907f
cc_44 N_Y_23 N_B_1 0.000783866f
cc_45 N_Y_19 N_MM1@2_g 0.0309692f
cc_46 N_Y_5 N_MM4@2_g 0.000890621f
cc_47 N_Y_2 N_B_8 0.0011574f
cc_48 N_Y_4 N_MM4@2_g 0.00222948f
cc_49 N_Y_17 N_MM1_g 0.0108225f
cc_50 N_Y_21 N_B_10 0.00563822f
cc_51 N_Y_19 N_B_1 0.006366f
cc_52 N_Y_20 N_MM4@2_g 0.0535019f
cc_53 N_Y_18 N_MM4@2_g 0.0212007f
cc_54 N_Y_19 N_MM1_g 0.0322022f
cc_55 N_Y_18 N_MM1@2_g 0.0503229f
cc_56 N_Y_3 N_NET16_15 0.00111967f
cc_57 N_Y_19 N_NET16_15 0.000556245f
cc_58 N_Y_20 N_NET16_15 0.00056063f
cc_59 N_Y_23 N_NET16_15 0.000642284f
cc_60 N_Y_22 N_NET16_3 0.000920998f
cc_61 N_Y_20 N_NET16_13 0.0011107f
cc_62 N_Y_19 N_NET16_13 0.00111424f
cc_63 N_Y_3 N_NET16_2 0.0011685f
cc_64 N_Y_3 N_NET16_3 0.00316164f
cc_65 N_Y_5 N_NET16_3 0.00432107f
cc_66 N_Y_22 N_NET16_15 0.0101703f
*END of NOR2x1p5_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR2x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR2x2_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00462958f
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0046437f
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00584743f
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00589499f
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%A VSS 29 3 4 5 6 7 1 8
c1 1 VSS 0.0209397f
c2 3 VSS 0.0843748f
c3 4 VSS 0.047223f
c4 5 VSS 0.0472272f
c5 6 VSS 0.0843454f
c6 7 VSS 0.00518702f
c7 8 VSS 0.00483705f
r1 8 31 2.31754 $w=1.6e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0720 $X2=0.2700 $Y2=0.0870
r2 6 27 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1355
r3 5 21 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1355
r4 29 7 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2700 $Y2=0.1095
r5 7 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1095 $X2=0.2700 $Y2=0.0870
r6 4 15 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1355
r7 25 27 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1355 $X2=0.3510 $Y2=0.1355
r8 24 25 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1355 $X2=0.3385 $Y2=0.1355
r9 22 24 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1355 $X2=0.3240 $Y2=0.1355
r10 21 22 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1355 $X2=0.3095 $Y2=0.1355
r11 19 21 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1355 $X2=0.2970 $Y2=0.1355
r12 18 19 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1355 $X2=0.2845 $Y2=0.1355
r13 29 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2700 $Y=0.1350
+ $X2=0.2700 $Y2=0.1355
r14 16 18 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1355 $X2=0.2700 $Y2=0.1355
r15 15 16 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1355 $X2=0.2555 $Y2=0.1355
r16 13 15 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1355 $X2=0.2430 $Y2=0.1355
r17 12 13 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1355 $X2=0.2305 $Y2=0.1355
r18 11 12 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1355 $X2=0.2160 $Y2=0.1355
r19 3 1 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1355
r20 1 10 2.59554 $w=2.2681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1355 $X2=0.1785 $Y2=0.1355
r21 1 11 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1355 $X2=0.2015 $Y2=0.1355
r22 3 10 0.54388 $w=2.16967e-07 $l=1.05119e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1355
r23 3 11 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1355
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%Y VSS 64 35 56 58 60 76 79 81 84 4 3 1 2 6 5 23
+ 22 19 27 28 26 25 24 29 21 20 33 31
c1 1 VSS 0.00766832f
c2 2 VSS 0.00289629f
c3 3 VSS 0.00755066f
c4 4 VSS 0.00770567f
c5 5 VSS 0.00770264f
c6 6 VSS 0.00290973f
c7 19 VSS 0.00346132f
c8 20 VSS 0.00347045f
c9 21 VSS 0.00346747f
c10 22 VSS 0.0034509f
c11 23 VSS 0.00211955f
c12 24 VSS 0.00211834f
c13 25 VSS 0.00227382f
c14 26 VSS 0.0392933f
c15 27 VSS 0.00064567f
c16 28 VSS 0.000698022f
c17 29 VSS 0.00237008f
c18 30 VSS 0.00283197f
c19 31 VSS 0.000792262f
c20 32 VSS 0.00298108f
c21 33 VSS 0.000792445f
r1 84 83 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 82 83 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 6 82 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.2025 $X2=0.4420 $Y2=0.2025
r4 24 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r5 81 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r6 79 78 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r7 2 78 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r8 75 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.2025 $X2=0.1100 $Y2=0.2025
r9 23 75 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.0980 $Y2=0.2025
r10 76 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r11 6 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r12 2 69 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r13 73 74 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r14 71 74 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r15 28 33 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5020 $Y=0.1980 $X2=0.5130 $Y2=0.1980
r16 28 71 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5020
+ $Y=0.1980 $X2=0.4840 $Y2=0.1980
r17 68 69 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r18 67 68 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1980 $X2=0.0855 $Y2=0.1980
r19 27 31 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0380 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r20 27 67 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0380
+ $Y=0.1980 $X2=0.0560 $Y2=0.1980
r21 33 66 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1980 $X2=0.5130 $Y2=0.1800
r22 31 54 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.1800
r23 65 66 5.07188 $w=1.3e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1582 $X2=0.5130 $Y2=0.1800
r24 64 65 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1450 $X2=0.5130 $Y2=0.1582
r25 64 63 6.12123 $w=1.3e-08 $l=2.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1450 $X2=0.5130 $Y2=0.1187
r26 62 63 7.40378 $w=1.3e-08 $l=3.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0870 $X2=0.5130 $Y2=0.1187
r27 61 62 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0720 $X2=0.5130 $Y2=0.0870
r28 29 32 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0540 $X2=0.5130 $Y2=0.0360
r29 29 61 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0540 $X2=0.5130 $Y2=0.0720
r30 22 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r31 60 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r32 58 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r33 21 57 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r34 20 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r35 56 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r36 53 54 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1260 $X2=0.0270 $Y2=0.1800
r37 52 53 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.1260
r38 25 30 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r39 25 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0720
r40 32 51 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.0360 $X2=0.4860 $Y2=0.0360
r41 5 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r42 4 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3275 $Y2=0.0360
r43 3 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2125 $Y2=0.0360
r44 30 37 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0540 $Y2=0.0360
r45 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r46 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4455
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r47 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r48 47 48 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r49 46 47 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3275
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r50 45 46 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3185
+ $Y=0.0360 $X2=0.3275 $Y2=0.0360
r51 44 45 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3185 $Y2=0.0360
r52 43 44 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2605
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r53 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.0360 $X2=0.2605 $Y2=0.0360
r54 41 42 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2215
+ $Y=0.0360 $X2=0.2335 $Y2=0.0360
r55 40 41 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2125
+ $Y=0.0360 $X2=0.2215 $Y2=0.0360
r56 39 40 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2125 $Y2=0.0360
r57 38 39 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1130
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r58 36 38 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1040
+ $Y=0.0360 $X2=0.1130 $Y2=0.0360
r59 26 36 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.0360 $X2=0.1040 $Y2=0.0360
r60 26 37 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r61 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1040 $Y2=0.0360
r62 35 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r63 19 34 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r64 4 21 1e-05
r65 1 19 1e-05
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%B VSS 35 5 6 7 8 12 1 2 10 18 14 20 17 13 11 19
+ 21 16 22 9 15
c1 1 VSS 0.00659001f
c2 2 VSS 0.00660597f
c3 5 VSS 0.00757101f
c4 6 VSS 0.0447944f
c5 7 VSS 0.0447977f
c6 8 VSS 0.00755915f
c7 9 VSS 0.00294257f
c8 10 VSS 0.00371414f
c9 11 VSS 0.00285025f
c10 12 VSS 0.00455035f
c11 13 VSS 0.0028551f
c12 14 VSS 0.00370556f
c13 15 VSS 0.00301248f
c14 16 VSS 0.00308043f
c15 17 VSS 0.00250446f
c16 18 VSS 0.00284437f
c17 19 VSS 0.00299752f
c18 20 VSS 0.00288841f
c19 21 VSS 0.00302634f
c20 22 VSS 0.00249651f
r1 7 55 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r2 8 48 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r3 53 55 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r4 52 53 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r5 50 52 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r6 2 48 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r7 2 50 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4465 $Y2=0.1350
r8 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1485
r9 46 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r10 15 46 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1095 $X2=0.4590 $Y2=0.1350
r11 22 45 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1620 $X2=0.4340 $Y2=0.1620
r12 22 47 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1620 $X2=0.4590 $Y2=0.1485
r13 14 20 9.45156 $w=1.34118e-08 $l=4.83141e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3790 $Y=0.1620 $X2=0.3310 $Y2=0.1675
r14 14 45 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3790
+ $Y=0.1620 $X2=0.4340 $Y2=0.1620
r15 13 21 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.1800 $X2=0.3310 $Y2=0.1980
r16 13 20 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3310 $Y=0.1800 $X2=0.3310 $Y2=0.1675
r17 21 43 5.46317 $w=1.44754e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3310 $Y=0.1980 $X2=0.3005 $Y2=0.1980
r18 42 43 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.3005 $Y2=0.1980
r19 41 42 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2515
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r20 12 19 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2300 $Y=0.1980 $X2=0.2090 $Y2=0.1980
r21 12 41 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2300
+ $Y=0.1980 $X2=0.2515 $Y2=0.1980
r22 11 40 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2090 $Y=0.1800 $X2=0.2090 $Y2=0.1675
r23 11 19 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.1800 $X2=0.2090 $Y2=0.1980
r24 18 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2090
+ $Y=0.1585 $X2=0.2090 $Y2=0.1675
r25 39 40 9.45156 $w=1.34118e-08 $l=4.83141e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1610 $Y=0.1620 $X2=0.2090 $Y2=0.1675
r26 38 39 10.6101 $w=1.3e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1155
+ $Y=0.1620 $X2=0.1610 $Y2=0.1620
r27 10 17 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0995 $Y=0.1620 $X2=0.0810 $Y2=0.1620
r28 10 38 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0995
+ $Y=0.1620 $X2=0.1155 $Y2=0.1620
r29 17 36 0.507892 $w=2.25351e-08 $l=9.3e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1620 $X2=0.0810 $Y2=0.1527
r30 35 36 0.174892 $w=1.3e-08 $l=7e-10 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1520 $X2=0.0810 $Y2=0.1527
r31 35 34 0.991057 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1520 $X2=0.0810 $Y2=0.1477
r32 33 34 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1477
r33 9 33 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1035 $X2=0.0810 $Y2=0.1350
r34 9 16 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1035 $X2=0.0810 $Y2=0.0720
r35 5 29 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r36 29 30 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r37 29 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r38 26 30 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.0905 $Y2=0.1350
r39 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r40 24 25 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r41 6 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r42 1 24 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r43 1 32 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1460 $Y2=0.1350
r44 6 24 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r45 6 32 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1460 $Y2=0.1350
.ends

.subckt PM_NOR2x2_ASAP7_75t_R%NET16 VSS 24 25 42 43 46 47 49 51 16 21 1 5 3 17
+ 20 19 4 2 18
c1 1 VSS 0.00524232f
c2 2 VSS 0.00708698f
c3 3 VSS 0.00909795f
c4 4 VSS 0.00724917f
c5 5 VSS 0.00525765f
c6 16 VSS 0.00221226f
c7 17 VSS 0.00332716f
c8 18 VSS 0.00435971f
c9 19 VSS 0.00333386f
c10 20 VSS 0.00221065f
c11 21 VSS 0.0386431f
r1 20 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 51 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 49 48 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r4 16 48 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r5 47 45 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r6 2 45 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r7 17 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r8 46 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r9 43 41 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r10 3 41 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r11 18 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r12 42 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r13 5 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r14 1 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r15 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r16 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r17 37 38 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r18 36 37 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4025
+ $Y=0.2340 $X2=0.4475 $Y2=0.2340
r19 35 36 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4025 $Y2=0.2340
r20 34 35 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3545
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r21 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0925 $Y2=0.2340
r22 29 30 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1855 $Y2=0.2340
r23 28 29 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1375
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r24 28 33 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1375
+ $Y=0.2340 $X2=0.0925 $Y2=0.2340
r25 27 34 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3095
+ $Y=0.2340 $X2=0.3545 $Y2=0.2340
r26 26 27 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3095 $Y2=0.2340
r27 21 26 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2305
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r28 21 30 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2305
+ $Y=0.2340 $X2=0.1855 $Y2=0.2340
r29 4 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r30 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r31 4 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r32 19 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r33 25 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r34 1 16 1e-05
.ends


*
.SUBCKT NOR2x2_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 VSS N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 VSS N_MM4@3_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@4 N_MM4@4_d N_MM1_g N_MM4@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM2_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@4 VDD N_MM3@4_g N_MM3@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@3 VDD N_MM3@3_g N_MM3@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 VDD N_MM2@2_g N_MM3@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM4@3_g N_MM4@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR2x2_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1 PM_NOR2x2_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM4_g 0.00920203f
cc_2 N_noxref_7_1 N_NET16_16 0.000639587f
cc_3 N_noxref_7_1 N_Y_19 0.00183301f
x_PM_NOR2x2_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_NOR2x2_ASAP7_75t_R%noxref_9
cc_4 N_noxref_9_1 N_MM4@2_g 0.0091512f
cc_5 N_noxref_9_1 N_NET16_20 0.000638397f
cc_6 N_noxref_9_1 N_Y_29 0.00047588f
cc_7 N_noxref_9_1 N_Y_22 0.0014033f
x_PM_NOR2x2_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1 PM_NOR2x2_ASAP7_75t_R%noxref_8
cc_8 N_noxref_8_1 N_MM4_g 0.00166587f
cc_9 N_noxref_8_1 N_NET16_16 0.0362085f
cc_10 N_noxref_8_1 N_Y_23 0.000791278f
cc_11 N_noxref_8_1 N_noxref_7_1 0.00193398f
x_PM_NOR2x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR2x2_ASAP7_75t_R%noxref_10
cc_12 N_noxref_10_1 N_MM4@2_g 0.001666f
cc_13 N_noxref_10_1 N_NET16_20 0.036157f
cc_14 N_noxref_10_1 N_Y_24 0.000790868f
cc_15 N_noxref_10_1 N_noxref_9_1 0.00193818f
x_PM_NOR2x2_ASAP7_75t_R%A VSS A N_MM2_g N_MM3@4_g N_MM3@3_g N_MM2@2_g N_A_7
+ N_A_1 N_A_8 PM_NOR2x2_ASAP7_75t_R%A
cc_16 N_MM2@2_g N_B_12 0.000276878f
cc_17 N_MM2@2_g N_B_1 0.000443022f
cc_18 N_MM2@2_g N_B_2 0.000444752f
cc_19 N_MM2@2_g N_B_10 0.00060935f
cc_20 N_MM2@2_g N_B_18 0.000611778f
cc_21 N_MM2@2_g N_B_14 0.000626726f
cc_22 N_A_7 N_B_12 0.00132999f
cc_23 N_A_1 N_B_12 0.00229684f
cc_24 N_A_7 N_B_20 0.0027246f
cc_25 N_MM2_g N_MM1_g 0.00337014f
cc_26 N_MM2@2_g N_MM4@3_g 0.00446955f
x_PM_NOR2x2_ASAP7_75t_R%Y VSS Y N_MM1_s N_MM2_s N_MM2@2_s N_MM1@2_s N_MM4_s
+ N_MM4@4_s N_MM4@3_s N_MM4@2_s N_Y_4 N_Y_3 N_Y_1 N_Y_2 N_Y_6 N_Y_5 N_Y_23
+ N_Y_22 N_Y_19 N_Y_27 N_Y_28 N_Y_26 N_Y_25 N_Y_24 N_Y_29 N_Y_21 N_Y_20 N_Y_33
+ N_Y_31 PM_NOR2x2_ASAP7_75t_R%Y
cc_27 N_Y_4 N_MM4@2_g 0.000273187f
cc_28 N_Y_3 N_B_18 0.000160546f
cc_29 N_Y_4 N_MM4@3_g 0.000177631f
cc_30 N_Y_3 N_MM1_g 0.000194795f
cc_31 N_Y_1 N_B_16 0.000340932f
cc_32 N_Y_2 N_B_10 0.0004243f
cc_33 N_Y_6 N_B_14 0.00044821f
cc_34 N_Y_1 N_B_1 0.00076686f
cc_35 N_Y_5 N_B_2 0.000882396f
cc_36 N_Y_23 N_MM1_g 0.0311155f
cc_37 N_Y_22 N_MM4@3_g 0.0492374f
cc_38 N_Y_19 N_MM1_g 0.070137f
cc_39 N_Y_6 N_MM4@2_g 0.00210337f
cc_40 N_Y_2 N_MM1_g 0.00210804f
cc_41 N_Y_27 N_B_10 0.00263196f
cc_42 N_Y_5 N_MM4@2_g 0.00263251f
cc_43 N_Y_28 N_B_14 0.0026458f
cc_44 N_Y_1 N_MM1_g 0.00293929f
cc_45 N_Y_26 N_B_16 0.00294401f
cc_46 N_Y_26 N_B_20 0.00389887f
cc_47 N_Y_28 N_B_22 0.0040174f
cc_48 N_Y_27 N_B_17 0.00430446f
cc_49 N_Y_23 N_B_1 0.00461448f
cc_50 N_Y_25 N_B_9 0.00463233f
cc_51 N_Y_24 N_B_2 0.00465815f
cc_52 N_Y_29 N_B_15 0.00489522f
cc_53 N_Y_22 N_MM4@2_g 0.0211763f
cc_54 N_Y_23 N_MM4_g 0.0378957f
cc_55 N_Y_24 N_MM4@2_g 0.0697388f
cc_56 N_Y_4 N_MM3@4_g 0.00110286f
cc_57 N_Y_21 N_MM3@4_g 0.0013024f
cc_58 N_Y_4 N_MM2@2_g 0.00256593f
cc_59 N_Y_3 N_MM3@4_g 0.00266643f
cc_60 N_Y_21 N_A_1 0.005142f
cc_61 N_Y_26 N_A_8 0.00582292f
cc_62 N_Y_21 N_MM3@3_g 0.0193229f
cc_63 N_Y_21 N_MM2@2_g 0.0503442f
cc_64 N_Y_20 N_MM2_g 0.0295274f
cc_65 N_Y_20 N_MM3@4_g 0.0426626f
cc_66 N_Y_2 N_NET16_21 0.000912389f
cc_67 N_Y_6 N_NET16_21 0.000988736f
cc_68 N_Y_27 N_NET16_1 0.000519904f
cc_69 N_Y_28 N_NET16_5 0.000519904f
cc_70 N_Y_24 N_NET16_19 0.000562395f
cc_71 N_Y_23 N_NET16_17 0.00168466f
cc_72 N_Y_33 N_NET16_21 0.000618717f
cc_73 N_Y_31 N_NET16_21 0.000626118f
cc_74 N_Y_23 N_NET16_16 0.000691481f
cc_75 N_Y_24 N_NET16_20 0.00181248f
cc_76 N_Y_29 N_NET16_5 0.000722044f
cc_77 N_Y_25 N_NET16_1 0.00073269f
cc_78 N_Y_6 N_NET16_4 0.00134079f
cc_79 N_Y_2 N_NET16_1 0.00238516f
cc_80 N_Y_27 N_NET16_21 0.00371426f
cc_81 N_Y_28 N_NET16_21 0.003726f
cc_82 N_Y_2 N_NET16_2 0.00409056f
cc_83 N_Y_6 N_NET16_5 0.00514662f
cc_84 N_Y_4 N_NET16_21 0.00877652f
x_PM_NOR2x2_ASAP7_75t_R%B VSS B N_MM4_g N_MM1_g N_MM4@3_g N_MM4@2_g N_B_12
+ N_B_1 N_B_2 N_B_10 N_B_18 N_B_14 N_B_20 N_B_17 N_B_13 N_B_11 N_B_19 N_B_21
+ N_B_16 N_B_22 N_B_9 N_B_15 PM_NOR2x2_ASAP7_75t_R%B
x_PM_NOR2x2_ASAP7_75t_R%NET16 VSS N_MM4@3_d N_MM3@2_s N_MM3@4_s N_MM3@3_s
+ N_MM4@4_d N_MM3_s N_MM4_d N_MM4@2_d N_NET16_16 N_NET16_21 N_NET16_1 N_NET16_5
+ N_NET16_3 N_NET16_17 N_NET16_20 N_NET16_19 N_NET16_4 N_NET16_2 N_NET16_18
+ PM_NOR2x2_ASAP7_75t_R%NET16
cc_85 N_NET16_16 N_B_17 0.000181705f
cc_86 N_NET16_21 N_B_13 0.000203646f
cc_87 N_NET16_21 N_B_11 0.000207906f
cc_88 N_NET16_1 N_B_1 0.000255424f
cc_89 N_NET16_5 N_B_2 0.00028906f
cc_90 N_NET16_3 N_B_12 0.00112208f
cc_91 N_NET16_17 N_MM1_g 0.0335084f
cc_92 N_NET16_20 N_MM4@2_g 0.0340419f
cc_93 N_NET16_19 N_MM4@3_g 0.0336168f
cc_94 N_NET16_21 N_B_19 0.00100857f
cc_95 N_NET16_21 N_B_21 0.00109293f
cc_96 N_NET16_1 N_MM4_g 0.00111979f
cc_97 N_NET16_5 N_MM4@2_g 0.0011207f
cc_98 N_NET16_4 N_B_14 0.00122255f
cc_99 N_NET16_2 N_B_10 0.00128239f
cc_100 N_NET16_4 N_MM4@3_g 0.00146579f
cc_101 N_NET16_2 N_MM1_g 0.00148655f
cc_102 N_NET16_20 N_B_2 0.00156306f
cc_103 N_NET16_17 N_B_1 0.00156987f
cc_104 N_NET16_21 N_B_12 0.0110507f
cc_105 N_NET16_16 N_MM4_g 0.0351915f
cc_106 N_NET16_17 N_MM3@3_g 0.000467413f
cc_107 N_NET16_4 N_MM3@3_g 0.000721617f
cc_108 N_NET16_2 N_MM3@3_g 0.000742052f
cc_109 N_NET16_3 N_MM3@3_g 0.00202448f
cc_110 N_NET16_18 N_A_1 0.00376312f
cc_111 N_NET16_19 N_MM2@2_g 0.0330496f
cc_112 N_NET16_17 N_MM2_g 0.0331493f
cc_113 N_NET16_18 N_MM3@4_g 0.0183837f
cc_114 N_NET16_18 N_MM3@3_g 0.0500787f
*END of NOR2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR2xp33_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR2xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR2xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR2xp33_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000842116f
r1 2 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r2 3 1 0.314815 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1080 $Y2=0.2160
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0317166f
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0208966f
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0205893f
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%A VSS 16 3 1 6 4 7
c1 1 VSS 0.00185125f
c2 3 VSS 0.04997f
c3 4 VSS 0.00508185f
c4 5 VSS 0.00541635f
c5 6 VSS 0.00138007f
c6 7 VSS 0.00710114f
c7 8 VSS 0.00108509f
c8 9 VSS 0.00767585f
r1 9 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 7 19 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r4 5 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r5 5 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r6 18 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 4 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 4 18 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 16 6 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 6 8 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r11 16 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r12 12 14 12.3648 $w=1.13e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r13 1 11 3.86521 $w=1.8e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r14 1 12 4.25053 $w=1.32143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r15 3 11 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r16 3 12 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00448626f
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%B VSS 4 3 1 5 6
c1 1 VSS 0.000862735f
c2 3 VSS 0.0220841f
c3 4 VSS 0.00445163f
c4 5 VSS 0.00174319f
c5 6 VSS 0.00345333f
r1 6 11 6.11415 $w=1.4371e-08 $l=3.1504e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1345 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 5 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 10 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r4 4 11 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1665
r5 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NOR2xp33_ASAP7_75t_R%Y VSS 23 16 17 28 7 9 1 8 11 2 10
c1 1 VSS 0.00671859f
c2 2 VSS 0.00600615f
c3 7 VSS 0.00354075f
c4 8 VSS 0.00301368f
c5 9 VSS 0.00899476f
c6 10 VSS 0.00396674f
c7 11 VSS 0.00477923f
c8 12 VSS 0.00362519f
c9 13 VSS 0.00302632f
r1 8 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1600 $Y2=0.2160
r2 28 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r3 2 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r4 10 13 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2340 $X2=0.1890 $Y2=0.2340
r5 13 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1890 $Y2=0.2160
r6 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.1890 $Y2=0.2160
r7 23 24 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1980
r8 23 22 14.691 $w=1.3e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0720
r9 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0360
r10 11 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0540 $X2=0.1890 $Y2=0.0720
r11 12 21 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0360 $X2=0.1620 $Y2=0.0360
r12 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1305
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r13 19 20 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r14 18 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1030
+ $Y=0.0360 $X2=0.1120 $Y2=0.0360
r15 9 18 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.0360 $X2=0.1030 $Y2=0.0360
r16 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0405
+ $X2=0.1120 $Y2=0.0360
r17 17 15 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0405 $X2=0.1225 $Y2=0.0405
r18 1 15 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0405 $X2=0.1225 $Y2=0.0405
r19 7 1 0.537037 $w=2.7e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0405 $X2=0.1080 $Y2=0.0405
r20 16 7 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0405 $X2=0.0935 $Y2=0.0405
.ends


*
.SUBCKT NOR2xp33_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM3 VDD N_MM2_g N_MM3_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NOR2xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR2xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR2xp33_ASAP7_75t_R%NET16 VSS N_MM3_s N_MM4_d N_NET16_1
+ PM_NOR2xp33_ASAP7_75t_R%NET16
cc_1 N_NET16_1 N_MM2_g 0.0125684f
cc_2 N_NET16_1 N_MM1_g 0.0125438f
x_PM_NOR2xp33_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NOR2xp33_ASAP7_75t_R%noxref_8
cc_3 N_noxref_8_1 N_MM2_g 0.004781f
cc_4 N_noxref_8_1 N_noxref_7_1 0.00202512f
x_PM_NOR2xp33_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NOR2xp33_ASAP7_75t_R%noxref_7
cc_5 N_noxref_7_1 N_MM2_g 0.00715045f
x_PM_NOR2xp33_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NOR2xp33_ASAP7_75t_R%noxref_9
cc_6 N_noxref_9_1 N_MM1_g 0.00592545f
cc_7 N_noxref_9_1 N_Y_7 0.00138929f
x_PM_NOR2xp33_ASAP7_75t_R%A VSS A N_MM2_g N_A_1 N_A_6 N_A_4 N_A_7
+ PM_NOR2xp33_ASAP7_75t_R%A
x_PM_NOR2xp33_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR2xp33_ASAP7_75t_R%noxref_10
cc_8 N_noxref_10_1 N_MM1_g 0.00372386f
cc_9 N_noxref_10_1 N_Y_8 0.0282188f
cc_10 N_noxref_10_1 N_noxref_9_1 0.00207849f
x_PM_NOR2xp33_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_5 N_B_6
+ PM_NOR2xp33_ASAP7_75t_R%B
cc_11 N_B_1 N_A_1 0.00266368f
cc_12 N_B_5 N_A_6 0.000555156f
cc_13 N_B_6 N_A_6 0.000659238f
cc_14 N_B N_A_6 0.00206852f
cc_15 N_MM1_g N_MM2_g 0.0122288f
x_PM_NOR2xp33_ASAP7_75t_R%Y VSS Y N_MM2_s N_MM1_s N_MM4_s N_Y_7 N_Y_9 N_Y_1
+ N_Y_8 N_Y_11 N_Y_2 N_Y_10 PM_NOR2xp33_ASAP7_75t_R%Y
cc_16 N_Y_7 N_A_6 0.000222078f
cc_17 N_Y_9 N_A_4 0.000280341f
cc_18 N_Y_1 N_MM2_g 0.000352475f
cc_19 N_Y_9 N_A_7 0.000864317f
cc_20 N_Y_7 N_MM2_g 0.0166268f
cc_21 N_Y_8 N_B_5 0.000375191f
cc_22 N_Y_1 N_MM1_g 0.000482215f
cc_23 N_Y_11 N_B_1 0.000505674f
cc_24 N_Y_8 N_B_1 0.000624555f
cc_25 N_Y_2 N_MM1_g 0.00110197f
cc_26 N_Y_7 N_MM1_g 0.00667028f
cc_27 N_Y_10 N_B_6 0.00259194f
cc_28 N_Y_9 N_B_5 0.00476261f
cc_29 N_Y_11 N_B 0.00628362f
cc_30 N_Y_8 N_MM1_g 0.0345093f
*END of NOR2xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR2xp67_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR2xp67_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR2xp67_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR2xp67_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00508722f
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00496005f
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0318821f
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00509173f
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%Y VSS 31 17 26 38 41 8 1 9 10 13 2 11 12 15
c1 1 VSS 0.0131743f
c2 2 VSS 0.00291694f
c3 8 VSS 0.0029405f
c4 9 VSS 0.00287034f
c5 10 VSS 0.00213492f
c6 11 VSS 0.0147275f
c7 12 VSS 0.000810553f
c8 13 VSS 0.00269832f
c9 14 VSS 0.00308401f
c10 15 VSS 0.000766119f
r1 41 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r2 39 40 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r3 2 39 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2160 $X2=0.2260 $Y2=0.2160
r4 10 2 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2140 $Y2=0.2160
r5 38 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r6 2 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.1980
r7 35 36 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2410 $Y2=0.1980
r8 33 36 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2705
+ $Y=0.1980 $X2=0.2410 $Y2=0.1980
r9 12 15 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2860 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r10 12 33 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2860
+ $Y=0.1980 $X2=0.2705 $Y2=0.1980
r11 15 32 3.30617 $w=1.71506e-08 $l=2.13e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1767
r12 31 32 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1640 $X2=0.2970 $Y2=0.1767
r13 31 30 2.39019 $w=1.3e-08 $l=1.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1640 $X2=0.2970 $Y2=0.1537
r14 29 30 4.37231 $w=1.3e-08 $l=1.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1537
r15 28 29 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1035 $X2=0.2970 $Y2=0.1350
r16 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.1035
r17 13 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0360
r18 13 27 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0720
r19 14 24 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2725 $Y2=0.0360
r20 26 25 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r21 9 25 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r22 23 24 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2140
+ $Y=0.0360 $X2=0.2725 $Y2=0.0360
r23 22 23 10.9599 $w=1.3e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1670
+ $Y=0.0360 $X2=0.2140 $Y2=0.0360
r24 21 22 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1580
+ $Y=0.0360 $X2=0.1670 $Y2=0.0360
r25 11 21 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1505
+ $Y=0.0360 $X2=0.1580 $Y2=0.0360
r26 9 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1580 $Y2=0.0360
r27 19 9 2.09809 $w=5.02e-08 $l=1.4e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1480 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r28 18 19 2.24795 $w=5.02e-08 $l=1.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1330 $Y=0.0540 $X2=0.1480 $Y2=0.0540
r29 1 18 3.74659 $w=5.02e-08 $l=2.5e-08 $layer=LISD $thickness=2.7e-08
+ $X=0.1080 $Y=0.0540 $X2=0.1330 $Y2=0.0540
r30 8 1 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1060 $Y2=0.0540
r31 17 8 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%B VSS 21 3 4 1 6 5 10 8 9 7
c1 1 VSS 0.00506657f
c2 3 VSS 0.0334791f
c3 4 VSS 0.0349251f
c4 5 VSS 0.00215235f
c5 6 VSS 0.00218232f
c6 7 VSS 0.00285097f
c7 8 VSS 0.00288211f
c8 9 VSS 0.00281198f
c9 10 VSS 0.00168258f
r1 8 26 6.04857 $w=1.44516e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1670
r2 6 25 0.983973 $w=1.77222e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1445 $X2=0.1350 $Y2=0.1355
r3 6 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1445 $X2=0.1350 $Y2=0.1670
r4 5 10 5.29779 $w=1.31087e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.1265
r5 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1035 $X2=0.1350 $Y2=0.0720
r6 10 24 2.26632 $w=1.325e-08 $l=2.03593e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1265 $X2=0.1535 $Y2=0.1350
r7 10 25 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1355
r8 23 24 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1825
+ $Y=0.1350 $X2=0.1535 $Y2=0.1350
r9 21 7 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2180 $Y2=0.1350
r10 7 23 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.1350 $X2=0.1825 $Y2=0.1350
r11 4 18 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1360
r12 21 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1360
r13 17 18 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1360 $X2=0.2430 $Y2=0.1360
r14 15 17 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1360 $X2=0.2335 $Y2=0.1360
r15 14 15 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1360 $X2=0.2305 $Y2=0.1360
r16 13 14 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1360 $X2=0.2160 $Y2=0.1360
r17 3 1 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1360
r18 1 12 3.05464 $w=2.15326e-08 $l=1.08e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1360 $X2=0.1782 $Y2=0.1360
r19 1 13 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1360 $X2=0.2015 $Y2=0.1360
r20 3 12 0.757708 $w=2.1223e-07 $l=1.08462e-08 $layer=LIG
+ $thickness=5.54419e-08 $X=0.1890 $Y=0.1350 $X2=0.1782 $Y2=0.1360
r21 3 13 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1360
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%NET16 VSS 15 28 31 33 1 2 10 13 11 3 12
c1 1 VSS 0.00698936f
c2 2 VSS 0.00589806f
c3 3 VSS 0.00510383f
c4 10 VSS 0.00322209f
c5 11 VSS 0.00292669f
c6 12 VSS 0.00221594f
c7 13 VSS 0.0203513f
r1 12 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2680 $Y2=0.2160
r2 33 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r3 31 30 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r4 2 30 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r5 27 2 0.222222 $w=5.4e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.2160 $X2=0.1640 $Y2=0.2160
r6 11 27 0.0833333 $w=5.4e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1520 $Y2=0.2160
r7 28 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r8 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r9 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r10 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r11 23 24 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1865
+ $Y=0.2340 $X2=0.2315 $Y2=0.2340
r12 22 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1865 $Y2=0.2340
r13 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r14 20 21 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1485 $Y2=0.2340
r15 19 20 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1010
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r16 18 19 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.2340 $X2=0.1010 $Y2=0.2340
r17 17 18 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0590
+ $Y=0.2340 $X2=0.0790 $Y2=0.2340
r18 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0500
+ $Y=0.2340 $X2=0.0590 $Y2=0.2340
r19 13 16 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0500 $Y2=0.2340
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0500 $Y2=0.2340
r21 15 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r22 10 14 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r23 1 10 1e-05
.ends

.subckt PM_NOR2xp67_ASAP7_75t_R%A VSS 22 3 4 1 7 10
c1 1 VSS 0.00294705f
c2 3 VSS 0.0593131f
c3 4 VSS 0.0317534f
c4 5 VSS 0.00849497f
c5 6 VSS 0.0038166f
c6 7 VSS 0.00202248f
c7 8 VSS 0.00889424f
c8 9 VSS 0.00193441f
c9 10 VSS 0.00347902f
r1 8 26 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 6 9 6.04857 $w=1.44516e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1670 $X2=0.0270 $Y2=0.1360
r3 6 10 6.04857 $w=1.44516e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1670 $X2=0.0270 $Y2=0.1980
r4 25 26 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r5 5 9 6.28176 $w=1.44063e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1040 $X2=0.0270 $Y2=0.1360
r6 5 25 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1040 $X2=0.0270 $Y2=0.0720
r7 9 24 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1360 $X2=0.0455 $Y2=0.1360
r8 4 20 2.92627 $w=1.245e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1360
r9 22 7 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0635 $Y2=0.1360
r10 7 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0635
+ $Y=0.1360 $X2=0.0455 $Y2=0.1360
r11 18 20 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1360 $X2=0.1350 $Y2=0.1360
r12 17 18 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1360 $X2=0.1225 $Y2=0.1360
r13 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1360 $X2=0.1080 $Y2=0.1360
r14 13 16 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1360 $X2=0.0935 $Y2=0.1360
r15 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0905 $Y2=0.1360
r16 22 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1360
+ $X2=0.0810 $Y2=0.1360
r17 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0810 $Y2=0.1360
r18 1 14 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0715 $Y=0.1360 $X2=0.0685 $Y2=0.1360
r19 3 12 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1360
r20 3 14 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1360
r21 3 16 1.79147 $w=1.8466e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1360
.ends


*
.SUBCKT NOR2xp67_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 VDD N_MM2_g N_MM3_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3@2 VDD N_MM3@2_g N_MM3@2_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2


*include "NOR2xp67_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR2xp67_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR2xp67_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NOR2xp67_ASAP7_75t_R%noxref_9
cc_1 N_noxref_9_1 N_MM4@2_g 0.00943815f
cc_2 N_noxref_9_1 N_NET16_12 0.000189219f
cc_3 N_noxref_9_1 N_Y_13 0.00140448f
x_PM_NOR2xp67_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR2xp67_ASAP7_75t_R%noxref_10
cc_4 N_noxref_10_1 N_MM4@2_g 0.00376f
cc_5 N_noxref_10_1 N_NET16_12 0.026794f
cc_6 N_noxref_10_1 N_Y_10 0.000954245f
cc_7 N_noxref_10_1 N_noxref_9_1 0.0021102f
x_PM_NOR2xp67_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_NOR2xp67_ASAP7_75t_R%noxref_7
cc_8 N_noxref_7_1 N_MM2_g 0.00471254f
x_PM_NOR2xp67_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_NOR2xp67_ASAP7_75t_R%noxref_8
cc_9 N_noxref_8_1 N_MM2_g 0.00463358f
cc_10 N_noxref_8_1 N_NET16_10 0.0268745f
cc_11 N_noxref_8_1 N_noxref_7_1 0.00203179f
x_PM_NOR2xp67_ASAP7_75t_R%Y VSS Y N_MM2_s N_MM1_s N_MM4_s N_MM4@2_s N_Y_8 N_Y_1
+ N_Y_9 N_Y_10 N_Y_13 N_Y_2 N_Y_11 N_Y_12 N_Y_15 PM_NOR2xp67_ASAP7_75t_R%Y
cc_12 N_Y_8 N_A_1 0.00101718f
cc_13 N_Y_1 N_MM3@2_g 0.00216265f
cc_14 N_Y_8 N_MM3@2_g 0.0147038f
cc_15 N_Y_8 N_MM2_g 0.0219205f
cc_16 N_Y_9 N_MM3@2_g 0.0417962f
cc_17 N_Y_1 N_MM1_g 0.000575179f
cc_18 N_Y_10 N_MM4@2_g 0.0363005f
cc_19 N_Y_13 N_B_1 0.00088795f
cc_20 N_Y_2 N_MM4@2_g 0.00090871f
cc_21 N_Y_10 N_B_1 0.00160679f
cc_22 N_Y_1 N_B_9 0.00168871f
cc_23 N_Y_13 N_B_7 0.00193736f
cc_24 N_Y_11 N_B_9 0.00434856f
cc_25 N_Y_12 N_B_7 0.00440413f
cc_26 N_Y_9 N_MM1_g 0.04015f
cc_27 N_Y_15 N_NET16_13 0.000607228f
cc_28 N_Y_12 N_NET16_3 0.000607246f
cc_29 N_Y_2 N_NET16_13 0.000742896f
cc_30 N_Y_10 N_NET16_12 0.000830601f
cc_31 N_Y_2 N_NET16_2 0.000998277f
cc_32 N_Y_2 N_NET16_3 0.0038809f
cc_33 N_Y_12 N_NET16_13 0.0101071f
x_PM_NOR2xp67_ASAP7_75t_R%B VSS B N_MM1_g N_MM4@2_g N_B_1 N_B_6 N_B_5 N_B_10
+ N_B_8 N_B_9 N_B_7 PM_NOR2xp67_ASAP7_75t_R%B
cc_34 N_B_1 N_A_1 0.000764855f
cc_35 N_B_6 N_A_7 0.000810842f
cc_36 N_B_5 N_A_7 0.000873603f
cc_37 N_B_10 N_A_7 0.00177883f
cc_38 N_B_10 N_A_1 0.00202164f
cc_39 N_MM1_g N_MM3@2_g 0.0102143f
x_PM_NOR2xp67_ASAP7_75t_R%NET16 VSS N_MM3_s N_MM3@2_s N_MM4_d N_MM4@2_d
+ N_NET16_1 N_NET16_2 N_NET16_10 N_NET16_13 N_NET16_11 N_NET16_3 N_NET16_12
+ PM_NOR2xp67_ASAP7_75t_R%NET16
cc_40 N_NET16_1 N_MM3@2_g 0.000449402f
cc_41 N_NET16_2 N_MM3@2_g 0.000452553f
cc_42 N_NET16_10 N_A_1 0.000719344f
cc_43 N_NET16_1 N_MM2_g 0.0012589f
cc_44 N_NET16_13 N_MM3@2_g 0.00155266f
cc_45 N_NET16_13 N_A_10 0.00184034f
cc_46 N_NET16_10 N_MM2_g 0.0242892f
cc_47 N_NET16_11 N_MM3@2_g 0.0258011f
cc_48 N_NET16_13 N_MM1_g 0.00050393f
cc_49 N_NET16_3 N_MM4@2_g 0.000537085f
cc_50 N_NET16_12 N_B_1 0.000595013f
cc_51 N_NET16_2 N_MM1_g 0.000839808f
cc_52 N_NET16_13 N_B_8 0.00539462f
cc_53 N_NET16_12 N_MM4@2_g 0.0241878f
cc_54 N_NET16_11 N_MM1_g 0.0259755f
x_PM_NOR2xp67_ASAP7_75t_R%A VSS A N_MM2_g N_MM3@2_g N_A_1 N_A_7 N_A_10
+ PM_NOR2xp67_ASAP7_75t_R%A
*END of NOR2xp67_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR3x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR3x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR3x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR3x1_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.00543446f
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0419623f
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%NET21 VSS 16 17 31 32 35 36 10 13 1 11 12 3 2
c1 1 VSS 0.00981597f
c2 2 VSS 0.00627262f
c3 3 VSS 0.00315393f
c4 10 VSS 0.00444709f
c5 11 VSS 0.00340855f
c6 12 VSS 0.00209858f
c7 13 VSS 0.0135223f
r1 36 34 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 34 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 35 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 32 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r6 2 30 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r8 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r9 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r10 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r11 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.1980 $X2=0.3240 $Y2=0.1980
r12 25 26 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2810
+ $Y=0.1980 $X2=0.3105 $Y2=0.1980
r13 24 25 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2450
+ $Y=0.1980 $X2=0.2810 $Y2=0.1980
r14 23 24 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.1980 $X2=0.2450 $Y2=0.1980
r15 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2295 $Y2=0.1980
r16 21 22 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r17 20 21 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.2045 $Y2=0.1980
r18 19 20 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r19 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1980 $X2=0.1465 $Y2=0.1980
r20 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.1980 $X2=0.1080 $Y2=0.1980
r21 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.1980
r22 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r23 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r24 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r25 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00531731f
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00468006f
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%B VSS 8 3 4 5 10 1 7 6 9
c1 1 VSS 0.0147133f
c2 3 VSS 0.04609f
c3 4 VSS 0.0481568f
c4 5 VSS 0.0483222f
c5 6 VSS 0.00575592f
c6 7 VSS 0.00445021f
c7 8 VSS 0.0053033f
c8 9 VSS 0.00451776f
c9 10 VSS 0.00389275f
r1 7 10 6.74572 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2610
+ $Y=0.1620 $X2=0.2970 $Y2=0.1620
r2 6 9 6.74572 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2610
+ $Y=0.0720 $X2=0.2970 $Y2=0.0720
r3 10 26 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1620 $X2=0.2970 $Y2=0.1485
r4 9 25 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.2970 $Y2=0.1035
r5 5 23 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 8 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r7 8 25 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1035
r8 8 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1485
r9 4 17 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 21 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r11 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r12 18 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r13 17 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r14 15 17 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r15 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r16 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r17 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r18 1 12 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r19 1 13 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r20 3 12 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r21 3 13 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%NET22 VSS 16 17 28 31 33 36 1 10 11 2 3 12 13
c1 1 VSS 0.00453217f
c2 2 VSS 0.00446305f
c3 3 VSS 0.00451247f
c4 10 VSS 0.00214777f
c5 11 VSS 0.00213405f
c6 12 VSS 0.0020982f
c7 13 VSS 0.0204611f
r1 36 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 34 35 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2800 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 1 34 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2680 $Y=0.2025 $X2=0.2800 $Y2=0.2025
r4 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r5 33 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r6 31 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r7 2 30 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3800 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r8 27 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3680 $Y=0.2025 $X2=0.3800 $Y2=0.2025
r9 11 27 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3680 $Y2=0.2025
r10 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r11 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r12 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r13 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r14 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r15 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r16 21 26 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r17 20 23 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r18 13 18 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r19 13 20 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.2340 $X2=0.4070 $Y2=0.2340
r20 3 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r22 3 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r23 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r24 16 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%C VSS 31 3 4 5 8 1
c1 1 VSS 0.0134605f
c2 3 VSS 0.0453225f
c3 4 VSS 0.0820861f
c4 5 VSS 0.0803725f
c5 6 VSS 0.0113491f
c6 7 VSS 0.00661374f
c7 8 VSS 0.00452471f
c8 9 VSS 0.00944876f
c9 10 VSS 0.00317867f
c10 11 VSS 0.00851908f
r1 11 37 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.1800
r2 9 35 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r3 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1620 $X2=0.0270 $Y2=0.1800
r4 7 10 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1485 $X2=0.0270 $Y2=0.1350
r5 7 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1485 $X2=0.0270 $Y2=0.1620
r6 34 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r7 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r8 6 34 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r9 10 33 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0455 $Y2=0.1350
r10 31 8 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1350 $X2=0.0580 $Y2=0.1350
r11 8 33 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0580
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r12 3 25 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 4 17 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r14 24 25 1.90543 $w=2e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.0850
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 23 24 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1350 $X2=0.0850 $Y2=0.1350
r16 31 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0700 $Y=0.1350
+ $X2=0.0750 $Y2=0.1350
r17 21 24 4.39635 $w=1.80294e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.0850 $Y2=0.1350
r18 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r19 18 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r20 17 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r21 15 17 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r22 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r23 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r24 5 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r25 1 13 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r26 1 30 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
r27 5 13 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r28 5 30 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%A VSS 23 3 4 5 1 8 9 7 10 6
c1 1 VSS 0.00929589f
c2 3 VSS 0.0463111f
c3 4 VSS 0.00888559f
c4 5 VSS 0.00978321f
c5 6 VSS 0.00507298f
c6 7 VSS 0.0047135f
c7 8 VSS 0.00427417f
c8 9 VSS 0.00399398f
c9 10 VSS 0.00376917f
r1 7 10 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.1620 $X2=0.4590 $Y2=0.1620
r2 6 9 6.74572 $w=1.425e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.4230
+ $Y=0.0720 $X2=0.4590 $Y2=0.0720
r3 10 24 1.49895 $w=1.95333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1620 $X2=0.4590 $Y2=0.1485
r4 5 21 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 3 15 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r6 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1485
r7 23 8 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1035
r8 8 9 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1035 $X2=0.4590 $Y2=0.0720
r9 19 21 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r10 18 19 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r11 17 18 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r12 13 15 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r13 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r14 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r15 4 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r16 23 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r17 4 11 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r18 4 17 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
.ends

.subckt PM_NOR3x1_ASAP7_75t_R%Y VSS 38 24 25 36 48 50 53 1 13 17 2 3 4 14 19 18
+ 15 16
c1 1 VSS 0.0110992f
c2 2 VSS 0.00761972f
c3 3 VSS 0.00290837f
c4 4 VSS 0.00410102f
c5 13 VSS 0.00476222f
c6 14 VSS 0.00345384f
c7 15 VSS 0.00213567f
c8 16 VSS 0.00232823f
c9 17 VSS 0.0336024f
c10 18 VSS 0.00193166f
c11 19 VSS 0.00270549f
c12 20 VSS 0.002564f
c13 21 VSS 0.00109119f
r1 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 51 52 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4420 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 3 51 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4300 $Y=0.2025 $X2=0.4420 $Y2=0.2025
r4 15 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r5 50 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r6 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5380 $Y2=0.2025
r7 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r8 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1980
r9 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.1980
r10 45 46 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r11 43 46 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4840
+ $Y=0.1980 $X2=0.4545 $Y2=0.1980
r12 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1980 $X2=0.5535 $Y2=0.1980
r13 18 41 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5155
+ $Y=0.1980 $X2=0.5400 $Y2=0.1980
r14 18 43 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5155
+ $Y=0.1980 $X2=0.4840 $Y2=0.1980
r15 21 40 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1980 $X2=0.5670 $Y2=0.1800
r16 21 42 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5535 $Y2=0.1980
r17 39 40 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1492 $X2=0.5670 $Y2=0.1800
r18 38 39 5.18847 $w=1.3e-08 $l=2.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1270 $X2=0.5670 $Y2=0.1492
r19 38 37 7.52037 $w=1.3e-08 $l=3.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1270 $X2=0.5670 $Y2=0.0947
r20 19 20 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0540 $X2=0.5670 $Y2=0.0360
r21 19 37 9.50248 $w=1.3e-08 $l=4.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0540 $X2=0.5670 $Y2=0.0947
r22 14 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r23 36 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r24 20 34 10.9431 $w=1.38333e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5130 $Y2=0.0360
r25 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r26 33 34 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4545
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r27 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4545 $Y2=0.0360
r28 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4095
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r29 30 31 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.0360 $X2=0.4095 $Y2=0.0360
r30 29 30 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.0360 $X2=0.3670 $Y2=0.0360
r31 28 29 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3220 $Y2=0.0360
r32 27 28 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r33 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r34 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2045
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r35 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r36 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r37 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r38 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r39 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends


*
.SUBCKT NOR3x1_ASAP7_75t_R VSS VDD C B A Y
*
* VSS VSS
* VDD VDD
* C C
* B B
* A A
* Y Y
*
*

MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@3 N_MM8@3_d N_MM8@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@3 N_MM10@3_d N_MM10@3_g N_MM10@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM10@2_g N_MM10@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM12_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@3 N_MM11@3_d N_MM11@3_g N_MM11@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g N_MM11@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR3x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR3x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR3x1_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_NOR3x1_ASAP7_75t_R%noxref_9
cc_1 N_noxref_9_1 N_MM8_g 0.0109336f
x_PM_NOR3x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR3x1_ASAP7_75t_R%noxref_10
cc_2 N_noxref_10_1 N_MM8_g 0.00251912f
cc_3 N_noxref_10_1 N_noxref_9_1 0.00193045f
x_PM_NOR3x1_ASAP7_75t_R%NET21 VSS N_MM8_d N_MM8@3_d N_MM8@2_d N_MM10_s
+ N_MM10@3_s N_MM10@2_s N_NET21_10 N_NET21_13 N_NET21_1 N_NET21_11 N_NET21_12
+ N_NET21_3 N_NET21_2 PM_NOR3x1_ASAP7_75t_R%NET21
cc_4 N_NET21_10 N_C_8 0.000588394f
cc_5 N_NET21_10 N_MM14_g 0.000683982f
cc_6 N_NET21_13 N_C_1 0.00134973f
cc_7 N_NET21_1 N_MM8@3_g 0.00179932f
cc_8 N_NET21_10 N_C_1 0.00324288f
cc_9 N_NET21_11 N_MM14_g 0.0325323f
cc_10 N_NET21_10 N_MM8_g 0.0180891f
cc_11 N_NET21_10 N_MM8@3_g 0.0496618f
cc_12 N_NET21_12 N_MM13_g 0.000864785f
cc_13 N_NET21_12 N_B_10 0.00116503f
cc_14 N_NET21_3 N_MM10@2_g 0.00186925f
cc_15 N_NET21_12 N_B_1 0.00287634f
cc_16 N_NET21_13 N_B_7 0.00649687f
cc_17 N_NET21_11 N_MM13_g 0.0325803f
cc_18 N_NET21_12 N_MM10@3_g 0.0181216f
cc_19 N_NET21_12 N_MM10@2_g 0.04964f
x_PM_NOR3x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NOR3x1_ASAP7_75t_R%noxref_12
cc_20 N_noxref_12_1 N_MM11@2_g 0.00165625f
cc_21 N_noxref_12_1 N_Y_16 0.0374117f
cc_22 N_noxref_12_1 N_noxref_11_1 0.00193668f
x_PM_NOR3x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NOR3x1_ASAP7_75t_R%noxref_11
cc_23 N_noxref_11_1 N_MM11@2_g 0.00943234f
cc_24 N_noxref_11_1 N_Y_16 0.00216719f
x_PM_NOR3x1_ASAP7_75t_R%B VSS B N_MM13_g N_MM10@3_g N_MM10@2_g N_B_10 N_B_1
+ N_B_7 N_B_6 N_B_9 PM_NOR3x1_ASAP7_75t_R%B
cc_25 N_MM13_g N_MM14_g 0.00498997f
x_PM_NOR3x1_ASAP7_75t_R%NET22 VSS N_MM11@3_s N_MM11@2_s N_MM10@2_d N_MM11_s
+ N_MM10_d N_MM10@3_d N_NET22_1 N_NET22_10 N_NET22_11 N_NET22_2 N_NET22_3
+ N_NET22_12 N_NET22_13 PM_NOR3x1_ASAP7_75t_R%NET22
cc_26 N_NET22_1 N_MM10@3_g 0.00195307f
cc_27 N_NET22_10 N_B_1 0.00269512f
cc_28 N_NET22_11 N_MM10@2_g 0.032729f
cc_29 N_NET22_10 N_MM13_g 0.0181061f
cc_30 N_NET22_10 N_MM10@3_g 0.0506842f
cc_31 N_NET22_2 N_MM12_g 0.000987043f
cc_32 N_NET22_3 N_MM11@2_g 0.00181283f
cc_33 N_NET22_12 N_A_1 0.00269356f
cc_34 N_NET22_11 N_MM12_g 0.03286f
cc_35 N_NET22_12 N_MM11@3_g 0.0181908f
cc_36 N_NET22_12 N_MM11@2_g 0.0504247f
cc_37 N_NET22_11 N_NET21_13 0.00110537f
cc_38 N_NET22_10 N_NET21_12 0.00111508f
cc_39 N_NET22_1 N_NET21_2 0.00122901f
cc_40 N_NET22_1 N_NET21_3 0.00299053f
cc_41 N_NET22_2 N_NET21_3 0.004153f
cc_42 N_NET22_13 N_NET21_13 0.012684f
x_PM_NOR3x1_ASAP7_75t_R%C VSS C N_MM8_g N_MM8@3_g N_MM14_g N_C_8 N_C_1
+ PM_NOR3x1_ASAP7_75t_R%C
x_PM_NOR3x1_ASAP7_75t_R%A VSS A N_MM12_g N_MM11@3_g N_MM11@2_g N_A_1 N_A_8
+ N_A_9 N_A_7 N_A_10 N_A_6 PM_NOR3x1_ASAP7_75t_R%A
cc_43 N_MM12_g N_MM10@2_g 0.00564468f
x_PM_NOR3x1_ASAP7_75t_R%Y VSS Y N_MM14_d N_MM13_d N_MM12_d N_MM11@2_d N_MM11_d
+ N_MM11@3_d N_Y_1 N_Y_13 N_Y_17 N_Y_2 N_Y_3 N_Y_4 N_Y_14 N_Y_19 N_Y_18 N_Y_15
+ N_Y_16 PM_NOR3x1_ASAP7_75t_R%Y
cc_44 N_Y_1 N_MM14_g 0.000797637f
cc_45 N_Y_13 N_C_1 0.000908755f
cc_46 N_Y_13 N_MM14_g 0.0344036f
cc_47 N_Y_17 N_MM13_g 0.000481634f
cc_48 N_Y_13 N_B_1 0.000914893f
cc_49 N_Y_1 N_MM13_g 0.00122728f
cc_50 N_Y_17 N_B_6 0.00246819f
cc_51 N_Y_17 N_B_9 0.00515598f
cc_52 N_Y_13 N_MM13_g 0.0349913f
cc_53 N_Y_2 N_MM11@3_g 0.00365014f
cc_54 N_Y_3 N_MM11@3_g 0.00250085f
cc_55 N_Y_4 N_MM11@2_g 0.000882011f
cc_56 N_Y_14 N_MM12_g 0.0492145f
cc_57 N_Y_19 N_A_1 0.00124643f
cc_58 N_Y_2 N_A_8 0.00130949f
cc_59 N_Y_17 N_A_9 0.00148124f
cc_60 N_Y_18 N_A_7 0.00220609f
cc_61 N_Y_18 N_A_10 0.00407831f
cc_62 N_Y_15 N_A_1 0.00590134f
cc_63 N_Y_17 N_A_6 0.00711303f
cc_64 N_Y_16 N_MM11@2_g 0.0347575f
cc_65 N_Y_14 N_MM11@3_g 0.0212053f
cc_66 N_Y_15 N_MM11@3_g 0.0697952f
cc_67 N_Y_16 N_NET22_13 0.000559788f
cc_68 N_Y_15 N_NET22_13 0.000562734f
cc_69 N_Y_3 N_NET22_13 0.000741771f
cc_70 N_Y_15 N_NET22_12 0.0011048f
cc_71 N_Y_16 N_NET22_12 0.0011233f
cc_72 N_Y_3 N_NET22_2 0.0013276f
cc_73 N_Y_3 N_NET22_3 0.00278391f
cc_74 N_Y_4 N_NET22_3 0.0043999f
cc_75 N_Y_18 N_NET22_13 0.0104866f
*END of NOR3x1_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR3x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR3x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR3x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR3x2_ASAP7_75t_R%NET21 VSS 28 29 53 54 57 58 61 62 65 66 69 70 24
+ 20 4 19 5 2 1 6 25 23 22 3 21
c1 1 VSS 0.00310229f
c2 2 VSS 0.00609206f
c3 3 VSS 0.0095355f
c4 4 VSS 0.00954862f
c5 5 VSS 0.00617847f
c6 6 VSS 0.00334639f
c7 19 VSS 0.00211826f
c8 20 VSS 0.00338809f
c9 21 VSS 0.00437253f
c10 22 VSS 0.00436574f
c11 23 VSS 0.00336444f
c12 24 VSS 0.00211473f
c13 25 VSS 0.0334004f
r1 70 68 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8270 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r2 6 68 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8100 $Y=0.2025 $X2=0.8245 $Y2=0.2025
r3 24 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.2025 $X2=0.8100 $Y2=0.2025
r4 69 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.2025 $X2=0.7955 $Y2=0.2025
r5 66 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r6 5 64 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.2025 $X2=0.7165 $Y2=0.2025
r7 23 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2025 $X2=0.7020 $Y2=0.2025
r8 65 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2025 $X2=0.6875 $Y2=0.2025
r9 62 60 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r10 4 60 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r11 22 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5940 $Y2=0.2025
r12 61 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r13 58 56 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r14 3 56 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r15 21 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r16 57 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r17 54 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r18 2 52 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r19 20 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r20 53 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r21 6 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.2025
+ $X2=0.8100 $Y2=0.1980
r22 5 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2025
+ $X2=0.7020 $Y2=0.1980
r23 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.1980
r24 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1980
r25 2 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r26 48 49 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7720
+ $Y=0.1980 $X2=0.8100 $Y2=0.1980
r27 47 48 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7425
+ $Y=0.1980 $X2=0.7720 $Y2=0.1980
r28 46 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7335
+ $Y=0.1980 $X2=0.7425 $Y2=0.1980
r29 45 46 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7180
+ $Y=0.1980 $X2=0.7335 $Y2=0.1980
r30 44 45 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.1980 $X2=0.7180 $Y2=0.1980
r31 43 44 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6775
+ $Y=0.1980 $X2=0.7020 $Y2=0.1980
r32 42 43 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.6325
+ $Y=0.1980 $X2=0.6775 $Y2=0.1980
r33 41 42 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.1980 $X2=0.6325 $Y2=0.1980
r34 40 41 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5750
+ $Y=0.1980 $X2=0.5940 $Y2=0.1980
r35 39 40 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.1980 $X2=0.5750 $Y2=0.1980
r36 38 39 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5210
+ $Y=0.1980 $X2=0.5560 $Y2=0.1980
r37 37 38 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1980 $X2=0.5210 $Y2=0.1980
r38 36 37 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4475
+ $Y=0.1980 $X2=0.4860 $Y2=0.1980
r39 35 36 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4025
+ $Y=0.1980 $X2=0.4475 $Y2=0.1980
r40 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.4025 $Y2=0.1980
r41 33 34 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3625
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r42 32 33 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1980 $X2=0.3625 $Y2=0.1980
r43 31 32 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3085
+ $Y=0.1980 $X2=0.3470 $Y2=0.1980
r44 30 31 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.3085 $Y2=0.1980
r45 25 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r46 1 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r47 28 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r48 1 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r49 19 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r50 29 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00535318f
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00533073f
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00468242f
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00468447f
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%B VSS 32 5 6 7 8 9 10 12 1 2 15 13 11 14
c1 1 VSS 0.0175799f
c2 2 VSS 0.0175048f
c3 5 VSS 0.0496523f
c4 6 VSS 0.0495782f
c5 7 VSS 0.0474897f
c6 8 VSS 0.0474171f
c7 9 VSS 0.0495782f
c8 10 VSS 0.0496439f
c9 11 VSS 0.00646957f
c10 12 VSS 0.0123019f
c11 13 VSS 0.0064149f
c12 14 VSS 0.00567558f
c13 15 VSS 0.00565883f
r1 10 56 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.8370
+ $Y=0.1350 $X2=0.8370 $Y2=0.1350
r2 9 50 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r3 8 42 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r4 54 56 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8245 $Y=0.1350 $X2=0.8370 $Y2=0.1350
r5 53 54 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.8100 $Y=0.1350 $X2=0.8245 $Y2=0.1350
r6 51 53 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7955 $Y=0.1350 $X2=0.8100 $Y2=0.1350
r7 50 51 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7955 $Y2=0.1350
r8 48 50 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1350 $X2=0.7830 $Y2=0.1350
r9 47 48 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1350 $X2=0.7705 $Y2=0.1350
r10 45 47 12.4546 $w=1.33e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7435 $Y=0.1350 $X2=0.7560 $Y2=0.1350
r11 44 45 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7410 $Y=0.1350 $X2=0.7435 $Y2=0.1350
r12 41 42 2.22301 $w=2e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.7320
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r13 41 44 4.21574 $w=1.85111e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7320 $Y=0.1350 $X2=0.7410 $Y2=0.1350
r14 2 41 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.7220
+ $Y=0.1350 $X2=0.7320 $Y2=0.1350
r15 38 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7340 $Y=0.1350
+ $X2=0.7320 $Y2=0.1350
r16 37 38 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.1160 $X2=0.7340 $Y2=0.1350
r17 13 15 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7340 $Y=0.0935 $X2=0.7340 $Y2=0.0720
r18 13 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7340
+ $Y=0.0935 $X2=0.7340 $Y2=0.1160
r19 15 36 19.1048 $w=1.35056e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7340 $Y=0.0720 $X2=0.6450 $Y2=0.0720
r20 35 36 20.7539 $w=1.3e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.0720 $X2=0.6450 $Y2=0.0720
r21 12 14 22.7192 $w=1.34306e-08 $l=1.045e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.4515 $Y=0.0720 $X2=0.3470 $Y2=0.0720
r22 12 35 24.3683 $w=1.3e-08 $l=1.045e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.4515 $Y=0.0720 $X2=0.5560 $Y2=0.0720
r23 14 34 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3470 $Y=0.0720 $X2=0.3470 $Y2=0.0935
r24 32 11 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1350 $X2=0.3470 $Y2=0.1160
r25 11 34 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3470
+ $Y=0.1160 $X2=0.3470 $Y2=0.0935
r26 7 29 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r27 5 20 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r28 27 29 2.38179 $w=2e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3485
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r29 32 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3470 $Y=0.1350
+ $X2=0.3485 $Y2=0.1350
r30 25 27 3.87634 $w=1.88833e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3395 $Y=0.1350 $X2=0.3485 $Y2=0.1350
r31 24 25 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3370 $Y=0.1350 $X2=0.3395 $Y2=0.1350
r32 23 24 12.9528 $w=1.33e-08 $l=1.3e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3370 $Y2=0.1350
r33 22 23 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r34 18 20 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r35 17 18 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r36 16 17 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r37 6 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r38 1 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r39 1 22 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r40 6 16 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r41 6 22 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%C VSS 45 3 4 5 6 7 8 9 1
c1 1 VSS 0.0326263f
c2 3 VSS 0.0848741f
c3 4 VSS 0.0866451f
c4 5 VSS 0.0494073f
c5 6 VSS 0.0493887f
c6 7 VSS 0.0866536f
c7 8 VSS 0.0848754f
c8 9 VSS 0.00624531f
r1 8 43 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r2 7 37 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r3 45 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5560
+ $Y=0.1350 $X2=0.5560 $Y2=0.1160
r4 6 31 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r5 5 22 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r6 4 16 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r7 41 43 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r8 40 41 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r9 38 40 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r10 37 38 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
r11 35 37 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6085 $Y=0.1350 $X2=0.6210 $Y2=0.1350
r12 34 35 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5940 $Y=0.1350 $X2=0.6085 $Y2=0.1350
r13 32 34 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5795 $Y=0.1350 $X2=0.5940 $Y2=0.1350
r14 30 31 1.90543 $w=2e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.5710
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r15 30 32 4.39635 $w=1.80294e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5710 $Y=0.1350 $X2=0.5795 $Y2=0.1350
r16 29 30 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.5610
+ $Y=0.1350 $X2=0.5710 $Y2=0.1350
r17 45 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5560 $Y=0.1350
+ $X2=0.5610 $Y2=0.1350
r18 27 29 3.76121 $w=1.74231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5610 $Y2=0.1350
r19 26 27 4.98184 $w=1.33e-08 $l=5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5495
+ $Y=0.1350 $X2=0.5545 $Y2=0.1350
r20 25 26 11.9564 $w=1.33e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5375 $Y=0.1350 $X2=0.5495 $Y2=0.1350
r21 23 25 11.9564 $w=1.33e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5375 $Y2=0.1350
r22 22 23 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r23 20 22 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r24 19 20 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r25 17 19 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r26 16 17 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r27 14 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r28 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r29 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r30 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r31 1 11 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r32 1 12 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r33 3 11 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r34 3 12 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%NET22 VSS 15 18 31 34 37 38 12 2 3 11 10 1 13
c1 1 VSS 0.00452766f
c2 2 VSS 0.00459721f
c3 3 VSS 0.00433548f
c4 10 VSS 0.00209679f
c5 11 VSS 0.00208798f
c6 12 VSS 0.00204307f
c7 13 VSS 0.0190931f
r1 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2025 $X2=0.9865 $Y2=0.2025
r2 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9720 $Y=0.2025 $X2=0.9865 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.2025 $X2=0.9720 $Y2=0.2025
r4 37 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2025 $X2=0.9575 $Y2=0.2025
r5 34 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8810 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r6 2 33 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8660 $Y=0.2025 $X2=0.8785 $Y2=0.2025
r7 30 2 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.8540 $Y=0.2025 $X2=0.8660 $Y2=0.2025
r8 11 30 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8495 $Y=0.2025 $X2=0.8540 $Y2=0.2025
r9 31 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.8470 $Y=0.2025 $X2=0.8495 $Y2=0.2025
r10 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9720 $Y=0.2025
+ $X2=0.9720 $Y2=0.2340
r11 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8640 $Y=0.2025
+ $X2=0.8605 $Y2=0.2340
r12 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9335
+ $Y=0.2340 $X2=0.9720 $Y2=0.2340
r13 26 27 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.9035
+ $Y=0.2340 $X2=0.9335 $Y2=0.2340
r14 25 26 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.2340 $X2=0.9035 $Y2=0.2340
r15 24 25 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.8790
+ $Y=0.2340 $X2=0.8940 $Y2=0.2340
r16 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.8695
+ $Y=0.2340 $X2=0.8790 $Y2=0.2340
r17 22 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.8605
+ $Y=0.2340 $X2=0.8695 $Y2=0.2340
r18 21 22 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.8395
+ $Y=0.2340 $X2=0.8605 $Y2=0.2340
r19 20 21 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7945
+ $Y=0.2340 $X2=0.8395 $Y2=0.2340
r20 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.2340 $X2=0.7945 $Y2=0.2340
r21 13 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7445
+ $Y=0.2340 $X2=0.7560 $Y2=0.2340
r22 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7560 $Y2=0.2340
r23 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r24 16 17 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7660 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r25 1 16 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7540 $Y=0.2025 $X2=0.7660 $Y2=0.2025
r26 10 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.2025 $X2=0.7540 $Y2=0.2025
r27 15 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.2025 $X2=0.7415 $Y2=0.2025
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%NET22__2 VSS 15 18 30 33 36 37 10 2 1 11 12 3 13
c1 1 VSS 0.00434496f
c2 2 VSS 0.00446951f
c3 3 VSS 0.00456548f
c4 10 VSS 0.00204803f
c5 11 VSS 0.00209579f
c6 12 VSS 0.00209921f
c7 13 VSS 0.0198989f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 1 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 36 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 33 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r6 31 32 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2260 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r7 2 31 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2140 $Y=0.2025 $X2=0.2260 $Y2=0.2025
r8 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r9 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r10 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r11 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2180 $Y2=0.2340
r12 27 28 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1465 $Y2=0.2340
r13 25 28 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1840
+ $Y=0.2340 $X2=0.1465 $Y2=0.2340
r14 23 24 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.2090 $Y2=0.2340
r15 23 25 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1995
+ $Y=0.2340 $X2=0.1840 $Y2=0.2340
r16 21 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.2340 $X2=0.2405 $Y2=0.2340
r17 21 24 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2180
+ $Y=0.2340 $X2=0.2090 $Y2=0.2340
r18 13 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r19 13 22 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.2405 $Y2=0.2340
r20 3 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r21 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r22 3 17 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r23 14 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3140 $Y=0.2025 $X2=0.3260 $Y2=0.2025
r24 12 14 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3140 $Y2=0.2025
r25 15 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%A VSS 39 5 6 7 8 9 10 14 13 1 2 11 12 15
c1 1 VSS 0.0026876f
c2 2 VSS 0.00264554f
c3 5 VSS 0.00614987f
c4 6 VSS 0.00524023f
c5 7 VSS 0.042722f
c6 8 VSS 0.0427119f
c7 9 VSS 0.00523826f
c8 10 VSS 0.00617432f
c9 11 VSS 0.00496721f
c10 12 VSS 0.00460051f
c11 13 VSS 0.00121297f
c12 14 VSS 0.00140976f
c13 15 VSS 0.0952099f
r1 10 59 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r2 9 53 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9450
+ $Y=0.1350 $X2=0.9450 $Y2=0.1350
r3 8 46 0.314665 $w=2.27e-07 $l=0 $layer=Gate_1 $thickness=5.6e-08 $X=0.8910
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r4 57 59 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9865 $Y=0.1350 $X2=0.9990 $Y2=0.1350
r5 56 57 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9720 $Y=0.1350 $X2=0.9865 $Y2=0.1350
r6 54 56 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9575 $Y=0.1350 $X2=0.9720 $Y2=0.1350
r7 53 54 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9575 $Y2=0.1350
r8 51 53 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9325 $Y=0.1350 $X2=0.9450 $Y2=0.1350
r9 50 51 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9180 $Y=0.1350 $X2=0.9325 $Y2=0.1350
r10 49 50 13.451 $w=1.33e-08 $l=1.35e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9045 $Y=0.1350 $X2=0.9180 $Y2=0.1350
r11 48 49 2.49092 $w=1.33e-08 $l=2.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.9020 $Y=0.1350 $X2=0.9045 $Y2=0.1350
r12 45 46 2.54058 $w=2e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.8930
+ $Y=0.1350 $X2=0.8910 $Y2=0.1350
r13 45 48 3.53695 $w=1.92556e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.8930 $Y=0.1350 $X2=0.9020 $Y2=0.1350
r14 2 45 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.8830
+ $Y=0.1350 $X2=0.8930 $Y2=0.1350
r15 39 14 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8940 $Y=0.0810 $X2=0.8940
+ $Y2=0.0720
r16 42 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.8940 $Y=0.1350
+ $X2=0.8930 $Y2=0.1350
r17 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.1080 $X2=0.8940 $Y2=0.1350
r18 12 41 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.8940
+ $Y=0.0855 $X2=0.8940 $Y2=0.1080
r19 39 12 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.8940 $Y=0.0810 $X2=0.8940
+ $Y2=0.0855
r20 12 14 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8940 $Y=0.0855 $X2=0.8940 $Y2=0.0720
r21 39 38 82.899 $w=1.3e-08 $l=3.555e-07 $layer=M2 $thickness=3.6e-08 $X=0.8940
+ $Y=0.0810 $X2=0.5385 $Y2=0.0810
r22 37 38 82.899 $w=1.3e-08 $l=3.555e-07 $layer=M2 $thickness=3.6e-08 $X=0.1830
+ $Y=0.0810 $X2=0.5385 $Y2=0.0810
r23 15 37 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1715
+ $Y=0.0810 $X2=0.1830 $Y2=0.0810
r24 13 37 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1830 $Y=0.0720 $X2=0.1830
+ $Y2=0.0810
r25 5 30 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r26 6 24 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r27 33 34 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1080 $X2=0.1830 $Y2=0.1350
r28 11 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.0855 $X2=0.1830 $Y2=0.1080
r29 11 13 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1830 $Y=0.0855 $X2=0.1830 $Y2=0.0720
r30 11 37 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1830 $Y=0.0855 $X2=0.1830
+ $Y2=0.0810
r31 28 30 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r32 27 28 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r33 25 27 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r34 24 25 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r35 22 24 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r36 21 22 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r37 20 21 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r38 19 32 1.60969 $w=1.91625e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1955 $Y=0.1350 $X2=0.1995 $Y2=0.1350
r39 1 19 3.17572 $w=2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.1855
+ $Y=0.1350 $X2=0.1955 $Y2=0.1350
r40 7 1 2.37889 $w=1.45455e-07 $l=3.5e-09 $layer=LIG $thickness=5.28485e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1855 $Y2=0.1350
r41 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1855 $Y=0.1350
+ $X2=0.1830 $Y2=0.1350
r42 7 20 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r43 7 32 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
.ends

.subckt PM_NOR3x2_ASAP7_75t_R%Y VSS 74 43 66 67 70 71 78 91 93 96 98 100 103 7
+ 3 2 6 34 29 32 1 8 31 33 37 25 28 36 35 30 27 4 5 26
c1 1 VSS 0.00413147f
c2 2 VSS 0.00765466f
c3 3 VSS 0.00292038f
c4 4 VSS 0.0100038f
c5 5 VSS 0.00978286f
c6 6 VSS 0.00777269f
c7 7 VSS 0.00291723f
c8 8 VSS 0.00412898f
c9 25 VSS 0.00347757f
c10 26 VSS 0.00472331f
c11 27 VSS 0.0047181f
c12 28 VSS 0.0034626f
c13 29 VSS 0.0023444f
c14 30 VSS 0.00217115f
c15 31 VSS 0.00217165f
c16 32 VSS 0.00233627f
c17 33 VSS 0.00283081f
c18 34 VSS 0.0890227f
c19 35 VSS 0.0021122f
c20 36 VSS 0.00220132f
c21 37 VSS 0.0028122f
c22 38 VSS 0.00275918f
c23 39 VSS 0.00107517f
c24 40 VSS 0.00275918f
c25 41 VSS 0.00107517f
r1 103 102 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9350 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r2 101 102 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9280 $Y=0.2025 $X2=0.9325 $Y2=0.2025
r3 7 101 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9160 $Y=0.2025 $X2=0.9280 $Y2=0.2025
r4 31 7 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.2025 $X2=0.9160 $Y2=0.2025
r5 100 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.2025 $X2=0.9035 $Y2=0.2025
r6 32 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.0115 $Y=0.2025 $X2=1.0240 $Y2=0.2025
r7 98 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=1.0090 $Y=0.2025 $X2=1.0115 $Y2=0.2025
r8 96 95 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r9 3 95 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r10 92 3 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1520 $Y=0.2025 $X2=0.1640 $Y2=0.2025
r11 30 92 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1520 $Y2=0.2025
r12 93 30 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r13 91 90 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r14 29 90 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r15 7 88 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.2025
+ $X2=0.9180 $Y2=0.1980
r16 8 85 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=1.0260 $Y=0.2025
+ $X2=1.0260 $Y2=0.1980
r17 3 82 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.1980
r18 1 79 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.1980
r19 88 89 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.1980 $X2=0.9565 $Y2=0.1980
r20 85 86 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.0260
+ $Y=0.1980 $X2=1.0395 $Y2=0.1980
r21 36 85 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=1.0015
+ $Y=0.1980 $X2=1.0260 $Y2=0.1980
r22 36 89 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.0015
+ $Y=0.1980 $X2=0.9565 $Y2=0.1980
r23 81 82 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r24 80 81 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0785
+ $Y=0.1980 $X2=0.1235 $Y2=0.1980
r25 79 80 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.1980 $X2=0.0785 $Y2=0.1980
r26 35 79 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.1980 $X2=0.0540 $Y2=0.1980
r27 35 39 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r28 41 76 3.59766 $w=1.692e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1980 $X2=1.0530 $Y2=0.1755
r29 41 86 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.1980 $X2=1.0395 $Y2=0.1980
r30 39 63 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r31 28 6 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9035 $Y=0.0675 $X2=0.9160 $Y2=0.0675
r32 78 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9010 $Y=0.0675 $X2=0.9035 $Y2=0.0675
r33 75 76 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1447 $X2=1.0530 $Y2=0.1755
r34 74 75 4.13912 $w=1.3e-08 $l=1.77e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1270 $X2=1.0530 $Y2=0.1447
r35 74 73 5.42166 $w=1.3e-08 $l=2.33e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1270 $X2=1.0530 $Y2=0.1037
r36 72 73 7.40378 $w=1.3e-08 $l=3.17e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0720 $X2=1.0530 $Y2=0.1037
r37 37 40 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0540 $X2=1.0530 $Y2=0.0360
r38 37 72 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0540 $X2=1.0530 $Y2=0.0720
r39 71 69 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r40 5 69 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r41 27 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r42 70 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r43 67 65 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r44 4 65 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r45 26 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r46 66 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r47 62 63 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1225 $X2=0.0270 $Y2=0.1765
r48 61 62 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.1225
r49 33 38 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r50 33 61 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0720
r51 6 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9180 $Y=0.0675
+ $X2=0.9180 $Y2=0.0360
r52 40 60 14.0912 $w=1.36667e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0360 $X2=0.9855 $Y2=0.0360
r53 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0675
+ $X2=0.7020 $Y2=0.0360
r54 4 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r55 59 60 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.9180
+ $Y=0.0360 $X2=0.9855 $Y2=0.0360
r56 58 59 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9065
+ $Y=0.0360 $X2=0.9180 $Y2=0.0360
r57 57 58 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.9035
+ $Y=0.0360 $X2=0.9065 $Y2=0.0360
r58 56 57 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.8845
+ $Y=0.0360 $X2=0.9035 $Y2=0.0360
r59 55 56 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.8450
+ $Y=0.0360 $X2=0.8845 $Y2=0.0360
r60 54 55 14.3412 $w=1.3e-08 $l=6.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7835
+ $Y=0.0360 $X2=0.8450 $Y2=0.0360
r61 53 54 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.7270
+ $Y=0.0360 $X2=0.7835 $Y2=0.0360
r62 52 53 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0360 $X2=0.7270 $Y2=0.0360
r63 51 52 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.7020 $Y2=0.0360
r64 50 51 37.7767 $w=1.3e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r65 49 50 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r66 48 49 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3535 $Y2=0.0360
r67 47 48 14.8076 $w=1.3e-08 $l=6.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2335
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r68 46 47 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1925
+ $Y=0.0360 $X2=0.2335 $Y2=0.0360
r69 45 46 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1725
+ $Y=0.0360 $X2=0.1925 $Y2=0.0360
r70 44 45 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1725 $Y2=0.0360
r71 34 44 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r72 34 38 14.0912 $w=1.36667e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r73 2 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r74 43 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r75 25 42 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1640 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r76 1 29 1e-05
r77 2 25 1e-05
.ends


*
.SUBCKT NOR3x2_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM10@5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM8_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14@2 N_MM14@2_d N_MM8@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13@2 N_MM13@2_d N_MM10_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12@2 N_MM12@2_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@4 N_MM11@4_d N_MM11@4_g N_MM11@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@6 N_MM11@6_d N_MM11@6_g N_MM11@6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@5 N_MM11@5_d N_MM12_g N_MM11@5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@4 N_MM10@4_d N_MM10@4_g N_MM10@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@6 N_MM10@6_d N_MM10@6_g N_MM10@6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@5 N_MM10@5_d N_MM10@5_g N_MM10@5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@6 N_MM8@6_d N_MM8@6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@5 N_MM8@5_d N_MM8@5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@4 N_MM8@4_d N_MM8@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@3 N_MM8@3_d N_MM8@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM8@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@3 N_MM10@3_d N_MM10@3_g N_MM10@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM10@2_g N_MM10@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@3 N_MM11@3_d N_MM11@3_g N_MM11@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g N_MM11@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR3x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR3x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR3x2_ASAP7_75t_R%NET21 VSS N_MM10@6_s N_MM10@4_s N_MM10@5_s N_MM8_d
+ N_MM8@6_d N_MM8@5_d N_MM8@4_d N_MM8@3_d N_MM8@2_d N_MM10_s N_MM10@3_s
+ N_MM10@2_s N_NET21_24 N_NET21_20 N_NET21_4 N_NET21_19 N_NET21_5 N_NET21_2
+ N_NET21_1 N_NET21_6 N_NET21_25 N_NET21_23 N_NET21_22 N_NET21_3 N_NET21_21
+ PM_NOR3x2_ASAP7_75t_R%NET21
cc_1 N_NET21_24 N_B_1 0.000351532f
cc_2 N_NET21_24 N_B_2 0.00345871f
cc_3 N_NET21_24 N_MM10_g 0.000427526f
cc_4 N_NET21_20 N_MM10@5_g 0.0330833f
cc_5 N_NET21_4 N_B_12 0.000755588f
cc_6 N_NET21_19 N_MM10@4_g 0.0480329f
cc_7 N_NET21_5 N_MM10_g 0.000884491f
cc_8 N_NET21_2 N_MM10@5_g 0.000890741f
cc_9 N_NET21_1 N_MM10@4_g 0.00164787f
cc_10 N_NET21_6 N_MM10@3_g 0.00165127f
cc_11 N_NET21_19 N_B_1 0.00313056f
cc_12 N_NET21_25 N_B_13 0.0036979f
cc_13 N_NET21_25 N_B_11 0.00380499f
cc_14 N_NET21_23 N_MM10_g 0.0325412f
cc_15 N_NET21_24 N_MM10@2_g 0.0180671f
cc_16 N_NET21_19 N_MM10@6_g 0.0181823f
cc_17 N_NET21_24 N_MM10@3_g 0.0489302f
cc_18 N_NET21_2 N_MM8@6_g 0.000673376f
cc_19 N_NET21_5 N_MM8@2_g 0.000683699f
cc_20 N_NET21_22 N_MM8@4_g 0.0482052f
cc_21 N_NET21_25 N_C_9 0.00165561f
cc_22 N_NET21_3 N_MM8@6_g 0.00168618f
cc_23 N_NET21_4 N_MM8@4_g 0.00173646f
cc_24 N_NET21_25 N_C_1 0.00241734f
cc_25 N_NET21_21 N_C_1 0.00635219f
cc_26 N_NET21_20 N_MM8_g 0.0325612f
cc_27 N_NET21_23 N_MM8@2_g 0.0326355f
cc_28 N_NET21_21 N_MM8@5_g 0.0181207f
cc_29 N_NET21_22 N_MM8@3_g 0.0181495f
cc_30 N_NET21_21 N_MM8@6_g 0.049844f
cc_31 N_NET21_1 N_NET22__2_13 0.000719995f
cc_32 N_NET21_19 N_NET22__2_11 0.00110863f
cc_33 N_NET21_19 N_NET22__2_12 0.00110879f
cc_34 N_NET21_2 N_NET22__2_3 0.00122538f
cc_35 N_NET21_1 N_NET22__2_3 0.00309836f
cc_36 N_NET21_1 N_NET22__2_2 0.00418956f
cc_37 N_NET21_25 N_NET22__2_13 0.0111143f
x_PM_NOR3x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NOR3x2_ASAP7_75t_R%noxref_11
cc_38 N_noxref_11_1 N_MM11@4_g 0.00166515f
cc_39 N_noxref_11_1 N_Y_33 0.000257134f
cc_40 N_noxref_11_1 N_Y_1 0.000493715f
cc_41 N_noxref_11_1 N_Y_29 0.0366625f
cc_42 N_noxref_11_1 N_noxref_10_1 0.00194147f
x_PM_NOR3x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NOR3x2_ASAP7_75t_R%noxref_13
cc_43 N_noxref_13_1 N_MM11@2_g 0.00166475f
cc_44 N_noxref_13_1 N_Y_37 0.000262262f
cc_45 N_noxref_13_1 N_Y_8 0.000493598f
cc_46 N_noxref_13_1 N_Y_32 0.0366822f
cc_47 N_noxref_13_1 N_noxref_12_1 0.00193959f
x_PM_NOR3x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR3x2_ASAP7_75t_R%noxref_10
cc_48 N_noxref_10_1 N_MM11@4_g 0.00943298f
cc_49 N_noxref_10_1 N_Y_34 0.000119481f
cc_50 N_noxref_10_1 N_Y_33 0.000512141f
cc_51 N_noxref_10_1 N_Y_29 0.00154659f
x_PM_NOR3x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NOR3x2_ASAP7_75t_R%noxref_12
cc_52 N_noxref_12_1 N_MM11@2_g 0.00941492f
cc_53 N_noxref_12_1 N_Y_34 0.000120016f
cc_54 N_noxref_12_1 N_Y_37 0.00051917f
cc_55 N_noxref_12_1 N_Y_32 0.00156357f
x_PM_NOR3x2_ASAP7_75t_R%B VSS B N_MM10@4_g N_MM10@6_g N_MM10@5_g N_MM10_g
+ N_MM10@3_g N_MM10@2_g N_B_12 N_B_1 N_B_2 N_B_15 N_B_13 N_B_11 N_B_14
+ PM_NOR3x2_ASAP7_75t_R%B
cc_56 N_B_12 N_A_14 8.9328e-20
cc_57 N_B_12 N_A_13 8.97689e-20
cc_58 N_B_12 N_A_1 9.78146e-20
cc_59 N_B_12 N_A_2 0.000108273f
cc_60 N_B_1 N_A_11 0.000219391f
cc_61 N_B_2 N_A_12 0.000229061f
cc_62 N_B_15 N_A_15 0.000317199f
cc_63 N_B_13 N_A_15 0.00106103f
cc_64 N_B_11 N_A_15 0.0011086f
cc_65 N_B_2 N_A_2 0.00115345f
cc_66 N_B_1 N_A_1 0.00117698f
cc_67 N_MM10@2_g N_MM11_g 0.00341735f
cc_68 N_MM10@4_g N_MM12_g 0.00341994f
cc_69 N_B_14 N_A_15 0.00389114f
cc_70 N_B_12 N_A_15 0.00847259f
x_PM_NOR3x2_ASAP7_75t_R%C VSS C N_MM8_g N_MM8@6_g N_MM8@5_g N_MM8@4_g N_MM8@3_g
+ N_MM8@2_g N_C_9 N_C_1 PM_NOR3x2_ASAP7_75t_R%C
cc_71 N_C_9 N_B_13 0.000173318f
cc_72 N_C_9 N_B_1 0.000352602f
cc_73 N_C_1 N_B_2 0.000355509f
cc_74 N_C_1 N_B_12 0.00266199f
cc_75 N_MM8@2_g N_MM10_g 0.00340201f
cc_76 N_MM8_g N_MM10@5_g 0.00340573f
cc_77 N_C_9 N_B_12 0.00663854f
x_PM_NOR3x2_ASAP7_75t_R%NET22 VSS N_MM10_d N_MM10@3_d N_MM10@2_d N_MM11_s
+ N_MM11@3_s N_MM11@2_s N_NET22_12 N_NET22_2 N_NET22_3 N_NET22_11 N_NET22_10
+ N_NET22_1 N_NET22_13 PM_NOR3x2_ASAP7_75t_R%NET22
cc_78 N_NET22_12 N_A_15 0.000288357f
cc_79 N_NET22_12 N_MM11_g 0.000419353f
cc_80 N_NET22_12 N_A_12 0.000983601f
cc_81 N_NET22_2 N_MM11_g 0.00103575f
cc_82 N_NET22_3 N_MM11@3_g 0.00164114f
cc_83 N_NET22_12 N_A_2 0.00268213f
cc_84 N_NET22_11 N_MM11_g 0.0326717f
cc_85 N_NET22_12 N_MM11@2_g 0.0180858f
cc_86 N_NET22_12 N_MM11@3_g 0.0483812f
cc_87 N_NET22_10 N_MM10@2_g 0.00114222f
cc_88 N_NET22_1 N_MM10_g 0.00180501f
cc_89 N_NET22_10 N_B_2 0.00277151f
cc_90 N_NET22_11 N_MM10@2_g 0.032553f
cc_91 N_NET22_10 N_MM10@3_g 0.0181542f
cc_92 N_NET22_10 N_MM10_g 0.0485581f
cc_93 N_NET22_13 N_NET21_6 0.000804942f
cc_94 N_NET22_10 N_NET21_24 0.00110937f
cc_95 N_NET22_10 N_NET21_23 0.00111001f
cc_96 N_NET22_2 N_NET21_6 0.00139686f
cc_97 N_NET22_1 N_NET21_6 0.00281538f
cc_98 N_NET22_1 N_NET21_5 0.00434741f
cc_99 N_NET22_13 N_NET21_25 0.01076f
x_PM_NOR3x2_ASAP7_75t_R%NET22__2 VSS N_MM10@6_d N_MM10@5_d N_MM11@5_s
+ N_MM10@4_d N_MM11@4_s N_MM11@6_s N_NET22__2_10 N_NET22__2_2 N_NET22__2_1
+ N_NET22__2_11 N_NET22__2_12 N_NET22__2_3 N_NET22__2_13
+ PM_NOR3x2_ASAP7_75t_R%NET22__2
cc_100 N_NET22__2_10 N_A_15 0.000298542f
cc_101 N_NET22__2_10 N_MM12_g 0.000450427f
cc_102 N_NET22__2_10 N_A_11 0.0010229f
cc_103 N_NET22__2_2 N_MM12_g 0.000999432f
cc_104 N_NET22__2_1 N_MM11@4_g 0.00165394f
cc_105 N_NET22__2_10 N_A_1 0.00268075f
cc_106 N_NET22__2_11 N_MM12_g 0.0327222f
cc_107 N_NET22__2_10 N_MM11@6_g 0.0181259f
cc_108 N_NET22__2_10 N_MM11@4_g 0.0484154f
cc_109 N_NET22__2_12 N_MM10@4_g 0.0011441f
cc_110 N_NET22__2_3 N_MM10@6_g 0.00183242f
cc_111 N_NET22__2_12 N_B_1 0.00280991f
cc_112 N_NET22__2_11 N_MM10@4_g 0.0326023f
cc_113 N_NET22__2_12 N_MM10@5_g 0.0180651f
cc_114 N_NET22__2_12 N_MM10@6_g 0.0487545f
x_PM_NOR3x2_ASAP7_75t_R%A VSS A N_MM11@4_g N_MM11@6_g N_MM12_g N_MM11_g
+ N_MM11@3_g N_MM11@2_g N_A_14 N_A_13 N_A_1 N_A_2 N_A_11 N_A_12 N_A_15
+ PM_NOR3x2_ASAP7_75t_R%A
x_PM_NOR3x2_ASAP7_75t_R%Y VSS Y N_MM12_d N_MM13_d N_MM14_d N_MM14@2_d
+ N_MM13@2_d N_MM12@2_d N_MM11@4_d N_MM11@6_d N_MM11@5_d N_MM11@2_d N_MM11_d
+ N_MM11@3_d N_Y_7 N_Y_3 N_Y_2 N_Y_6 N_Y_34 N_Y_29 N_Y_32 N_Y_1 N_Y_8 N_Y_31
+ N_Y_33 N_Y_37 N_Y_25 N_Y_28 N_Y_36 N_Y_35 N_Y_30 N_Y_27 N_Y_4 N_Y_5 N_Y_26
+ PM_NOR3x2_ASAP7_75t_R%Y
cc_115 N_Y_7 N_A_12 0.000252768f
cc_116 N_Y_3 N_A_11 0.000270477f
cc_117 N_Y_2 N_A_13 0.000331008f
cc_118 N_Y_6 N_A_14 0.000331171f
cc_119 N_Y_34 N_A_12 0.000344024f
cc_120 N_Y_34 N_A_11 0.000361574f
cc_121 N_Y_29 N_MM11@4_g 0.0352978f
cc_122 N_Y_32 N_MM11@2_g 0.0353146f
cc_123 N_Y_3 N_A_1 0.000596541f
cc_124 N_Y_7 N_A_2 0.000609166f
cc_125 N_Y_1 N_MM11@4_g 0.000838142f
cc_126 N_Y_8 N_MM11@2_g 0.000840446f
cc_127 N_Y_31 N_MM11_g 0.0309367f
cc_128 N_Y_33 N_A_1 0.00104354f
cc_129 N_Y_37 N_A_2 0.00107367f
cc_130 N_Y_25 N_MM12_g 0.0492255f
cc_131 N_Y_28 N_MM11_g 0.0703258f
cc_132 N_Y_36 N_A_2 0.00142197f
cc_133 N_Y_35 N_A_1 0.00152647f
cc_134 N_Y_6 N_A_12 0.00179911f
cc_135 N_Y_3 N_MM11@6_g 0.0018858f
cc_136 N_Y_7 N_MM11_g 0.00188657f
cc_137 N_Y_2 N_A_11 0.00202372f
cc_138 N_Y_34 N_A_13 0.00262864f
cc_139 N_Y_34 N_A_14 0.00271254f
cc_140 N_Y_6 N_MM11_g 0.00288343f
cc_141 N_Y_2 N_MM11@6_g 0.00293312f
cc_142 N_Y_30 N_A_1 0.00633061f
cc_143 N_Y_31 N_A_2 0.00641139f
cc_144 N_Y_34 N_A_15 0.0171256f
cc_145 N_Y_25 N_MM11@6_g 0.0211839f
cc_146 N_Y_31 N_MM11@3_g 0.0378309f
cc_147 N_Y_30 N_MM11@6_g 0.0691347f
cc_148 N_Y_27 N_MM10@5_g 0.000123597f
cc_149 N_Y_28 N_MM10@5_g 0.00014816f
cc_150 N_Y_25 N_MM10@5_g 0.000154083f
cc_151 N_Y_4 N_B_1 0.000184722f
cc_152 N_Y_5 N_B_2 0.000190845f
cc_153 N_Y_4 N_B_12 0.000426622f
cc_154 N_Y_27 N_MM10_g 0.0339843f
cc_155 N_Y_5 N_B_12 0.000449336f
cc_156 N_Y_5 N_B_13 0.000566709f
cc_157 N_Y_4 N_B_11 0.000596903f
cc_158 N_Y_26 N_B_1 0.000887916f
cc_159 N_Y_27 N_B_2 0.000957791f
cc_160 N_Y_4 N_MM10@5_g 0.00171095f
cc_161 N_Y_5 N_MM10_g 0.00174027f
cc_162 N_Y_34 N_B_15 0.0085401f
cc_163 N_Y_34 N_B_14 0.00877035f
cc_164 N_Y_34 N_B_12 0.0136872f
cc_165 N_Y_26 N_MM10@5_g 0.0344643f
cc_166 N_Y_26 N_MM8@2_g 0.00059083f
cc_167 N_Y_34 N_MM8@2_g 0.000593982f
cc_168 N_Y_4 N_MM8_g 0.000696063f
cc_169 N_Y_5 N_MM8@2_g 0.000731429f
cc_170 N_Y_34 N_C_1 0.00149254f
cc_171 N_Y_26 N_MM8_g 0.0335346f
cc_172 N_Y_27 N_MM8@2_g 0.0345315f
cc_173 N_Y_33 N_NET22__2_13 0.000137094f
cc_174 N_Y_1 N_NET22__2_13 0.000202076f
cc_175 N_Y_3 N_NET22__2_13 0.000957144f
cc_176 N_Y_30 N_NET22__2_13 0.0005562f
cc_177 N_Y_29 N_NET22__2_13 0.000556796f
cc_178 N_Y_30 N_NET22__2_10 0.00110975f
cc_179 N_Y_29 N_NET22__2_10 0.00112075f
cc_180 N_Y_3 N_NET22__2_2 0.00133504f
cc_181 N_Y_3 N_NET22__2_1 0.00277702f
cc_182 N_Y_1 N_NET22__2_1 0.00454861f
cc_183 N_Y_35 N_NET22__2_13 0.00944555f
cc_184 N_Y_37 N_NET22_13 0.000128804f
cc_185 N_Y_7 N_NET22_13 0.000955501f
cc_186 N_Y_8 N_NET22_13 0.000261443f
cc_187 N_Y_32 N_NET22_13 0.000554196f
cc_188 N_Y_31 N_NET22_13 0.000554413f
cc_189 N_Y_31 N_NET22_11 0.00110908f
cc_190 N_Y_31 N_NET22_12 0.00111793f
cc_191 N_Y_8 N_NET22_3 0.00126235f
cc_192 N_Y_7 N_NET22_3 0.00327716f
cc_193 N_Y_7 N_NET22_2 0.00412757f
cc_194 N_Y_36 N_NET22_13 0.00942805f
*END of NOR3x2_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR3xp33_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR3xp33_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR3xp33_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR3xp33_ASAP7_75t_R%NET22 VSS 2 3 1
c1 1 VSS 0.000896666f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%NET21 VSS 2 3 1
c1 1 VSS 0.000901044f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0425192f
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0327927f
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00379514f
c2 3 VSS 0.0716089f
c3 4 VSS 0.0159034f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0044025f
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00453968f
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00501188f
c2 3 VSS 0.0345851f
c3 4 VSS 0.00430121f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00430924f
c2 3 VSS 0.0354261f
c3 4 VSS 0.00709997f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NOR3xp33_ASAP7_75t_R%Y VSS 29 18 34 35 40 12 2 14 10 13 3 11
c1 2 VSS 0.00595084f
c2 3 VSS 0.00851998f
c3 10 VSS 0.00997417f
c4 11 VSS 0.00403134f
c5 12 VSS 0.00259297f
c6 13 VSS 0.00286013f
c7 14 VSS 0.0135539f
c8 15 VSS 0.00309027f
c9 16 VSS 0.00598355f
r1 40 39 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 12 39 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 16 31 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 16 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 35 33 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r8 3 33 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r9 11 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r10 34 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r11 30 31 11.368 $w=1.3e-08 $l=4.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1637 $X2=0.0270 $Y2=0.2125
r12 29 30 8.56972 $w=1.3e-08 $l=3.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1270 $X2=0.0270 $Y2=0.1637
r13 29 28 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1270 $X2=0.0270 $Y2=0.0982
r14 13 15 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r15 13 28 9.50248 $w=1.3e-08 $l=4.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.0982
r16 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r17 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r18 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1485 $Y2=0.0360
r19 23 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r20 22 23 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r21 21 22 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r22 20 21 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0655
+ $Y=0.0360 $X2=0.0700 $Y2=0.0360
r23 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0655 $Y2=0.0360
r24 14 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r25 14 15 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r26 10 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0000 $Y=0.0000
+ $X2=0.0540 $Y2=0.0360
r27 18 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r28 10 17 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r29 2 12 1e-05
.ends


*
.SUBCKT NOR3xp33_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM11 N_MM11_d N_MM12_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR3xp33_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR3xp33_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR3xp33_ASAP7_75t_R%NET22 VSS N_MM11_s N_MM10_d N_NET22_1
+ PM_NOR3xp33_ASAP7_75t_R%NET22
cc_1 N_NET22_1 N_MM12_g 0.0171874f
cc_2 N_NET22_1 N_MM13_g 0.0173121f
x_PM_NOR3xp33_ASAP7_75t_R%NET21 VSS N_MM10_s N_MM8_d N_NET21_1
+ PM_NOR3xp33_ASAP7_75t_R%NET21
cc_3 N_NET21_1 N_MM13_g 0.0172442f
cc_4 N_NET21_1 N_MM14_g 0.0172499f
x_PM_NOR3xp33_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NOR3xp33_ASAP7_75t_R%noxref_12
cc_5 N_noxref_12_1 N_MM14_g 0.0018487f
cc_6 N_noxref_12_1 N_noxref_11_1 0.0019265f
x_PM_NOR3xp33_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NOR3xp33_ASAP7_75t_R%noxref_11
cc_7 N_noxref_11_1 N_MM14_g 0.00377313f
x_PM_NOR3xp33_ASAP7_75t_R%C VSS C N_MM14_g N_C_1 N_C_4 PM_NOR3xp33_ASAP7_75t_R%C
cc_8 N_C_1 N_B_1 0.00159594f
cc_9 N_C_4 N_B_4 0.00669955f
cc_10 N_MM14_g N_MM13_g 0.00851086f
x_PM_NOR3xp33_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1
+ PM_NOR3xp33_ASAP7_75t_R%noxref_9
cc_11 N_noxref_9_1 N_MM12_g 0.0034879f
cc_12 N_noxref_9_1 N_Y_10 0.0288151f
x_PM_NOR3xp33_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_NOR3xp33_ASAP7_75t_R%noxref_10
cc_13 N_noxref_10_1 N_MM12_g 0.00160149f
cc_14 N_noxref_10_1 N_Y_12 0.0383568f
cc_15 N_noxref_10_1 N_noxref_9_1 0.00189375f
x_PM_NOR3xp33_ASAP7_75t_R%A VSS A N_MM12_g N_A_1 N_A_4 PM_NOR3xp33_ASAP7_75t_R%A
x_PM_NOR3xp33_ASAP7_75t_R%B VSS B N_MM13_g N_B_1 N_B_4 PM_NOR3xp33_ASAP7_75t_R%B
cc_16 N_B_1 N_A_1 0.00159238f
cc_17 N_B_4 N_A_4 0.00546137f
cc_18 N_MM13_g N_MM12_g 0.00843815f
x_PM_NOR3xp33_ASAP7_75t_R%Y VSS Y N_MM12_d N_MM13_d N_MM14_d N_MM11_d N_Y_12
+ N_Y_2 N_Y_14 N_Y_10 N_Y_13 N_Y_3 N_Y_11 PM_NOR3xp33_ASAP7_75t_R%Y
cc_19 N_Y_12 N_A_4 0.000489364f
cc_20 N_Y_2 N_A_1 0.000780318f
cc_21 N_Y_14 N_A_4 0.00108034f
cc_22 N_Y_12 N_A_1 0.00132423f
cc_23 N_Y_2 N_MM12_g 0.00171049f
cc_24 N_Y_10 N_MM12_g 0.0107419f
cc_25 N_Y_13 N_A_4 0.00787682f
cc_26 N_Y_12 N_MM12_g 0.0509328f
cc_27 N_Y_3 N_MM13_g 0.000607261f
cc_28 N_Y_14 N_B_4 0.00110513f
cc_29 N_Y_2 N_B_4 0.0020412f
cc_30 N_Y_11 N_MM13_g 0.0268853f
cc_31 N_Y_11 N_C_4 0.000601981f
cc_32 N_Y_3 N_C_4 0.00120982f
cc_33 N_Y_11 N_MM14_g 0.0263833f
*END of NOR3xp33_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR4xp25_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR4xp25_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR4xp25_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR4xp25_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0425498f
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%PD3 VSS 2 3 1
c1 1 VSS 0.000904734f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%PD1 VSS 2 3 1
c1 1 VSS 0.000893243f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%PD2 VSS 2 3 1
c1 1 VSS 0.000835994f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00497972f
c2 3 VSS 0.0345566f
c3 4 VSS 0.00428577f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00532631f
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00495868f
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.004524f
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%D VSS 10 3 1 4
c1 1 VSS 0.0036679f
c2 3 VSS 0.0714432f
c3 4 VSS 0.0150701f
r1 10 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 7 9 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1350 $X2=0.0915 $Y2=0.1350
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r4 10 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r6 1 8 2.51167 $w=1.2975e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0695 $Y2=0.1350
r7 3 6 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r8 3 8 2.63307 $w=1.98865e-07 $l=1.15e-08 $layer=LIG $thickness=5.49565e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0695 $Y2=0.1350
r9 3 9 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1350
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00435363f
c2 3 VSS 0.0356635f
c3 4 VSS 0.00741508f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00384476f
c2 3 VSS 0.0350368f
c3 4 VSS 0.00699177f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_NOR4xp25_ASAP7_75t_R%Y VSS 43 22 40 41 47 52 1 17 13 2 14 4 19 3 16
+ 15 18
c1 1 VSS 0.00759727f
c2 2 VSS 0.00839967f
c3 3 VSS 0.00681979f
c4 4 VSS 0.00614139f
c5 13 VSS 0.00338638f
c6 14 VSS 0.00391235f
c7 15 VSS 0.0031453f
c8 16 VSS 0.0025808f
c9 17 VSS 0.0231432f
c10 18 VSS 0.00289692f
c11 19 VSS 0.00594436f
c12 20 VSS 0.00306152f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 52 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 4 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r4 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r5 19 45 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2970 $Y2=0.2125
r6 19 50 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2835 $Y2=0.2340
r7 15 3 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0540 $X2=0.2680 $Y2=0.0540
r8 47 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2555 $Y2=0.0540
r9 44 45 11.7178 $w=1.3e-08 $l=5.03e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1622 $X2=0.2970 $Y2=0.2125
r10 43 44 8.91951 $w=1.3e-08 $l=3.82e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1240 $X2=0.2970 $Y2=0.1622
r11 43 42 6.35442 $w=1.3e-08 $l=2.73e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1240 $X2=0.2970 $Y2=0.0967
r12 18 20 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0575 $X2=0.2970 $Y2=0.0360
r13 18 42 9.1527 $w=1.3e-08 $l=3.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0575 $X2=0.2970 $Y2=0.0967
r14 41 39 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r15 2 39 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r16 14 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r17 40 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r18 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r19 20 37 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2835 $Y2=0.0360
r20 2 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r21 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r22 35 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r23 34 35 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2540
+ $Y=0.0360 $X2=0.2585 $Y2=0.0360
r24 33 34 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2540 $Y2=0.0360
r25 32 33 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r26 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r27 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r28 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r29 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r30 27 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1485 $Y2=0.0360
r31 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r32 25 26 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r33 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r34 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r35 17 23 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r36 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r37 22 21 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r38 13 21 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r39 1 13 1e-05
.ends


*
.SUBCKT NOR4xp25_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM1_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM0_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR4xp25_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR4xp25_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR4xp25_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NOR4xp25_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM3_g 0.00185757f
cc_2 N_noxref_12_1 N_noxref_11_1 0.00192378f
x_PM_NOR4xp25_ASAP7_75t_R%PD3 VSS N_MM4_d N_MM5_s N_PD3_1
+ PM_NOR4xp25_ASAP7_75t_R%PD3
cc_3 N_PD3_1 N_MM3_g 0.0172283f
cc_4 N_PD3_1 N_MM2_g 0.0173833f
x_PM_NOR4xp25_ASAP7_75t_R%PD1 VSS N_MM6_d N_MM7_s N_PD1_1
+ PM_NOR4xp25_ASAP7_75t_R%PD1
cc_5 N_PD1_1 N_MM1_g 0.0173348f
cc_6 N_PD1_1 N_MM0_g 0.0173963f
x_PM_NOR4xp25_ASAP7_75t_R%PD2 VSS N_MM5_d N_MM6_s N_PD2_1
+ PM_NOR4xp25_ASAP7_75t_R%PD2
cc_7 N_PD2_1 N_MM2_g 0.0172913f
cc_8 N_PD2_1 N_MM1_g 0.0173602f
x_PM_NOR4xp25_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_NOR4xp25_ASAP7_75t_R%A
cc_9 N_A_1 N_B_1 0.00151116f
cc_10 N_A_4 N_B_4 0.00548571f
cc_11 N_MM0_g N_MM1_g 0.00837153f
x_PM_NOR4xp25_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NOR4xp25_ASAP7_75t_R%noxref_11
cc_12 N_noxref_11_1 N_MM3_g 0.00373598f
cc_13 N_noxref_11_1 N_Y_13 0.0274367f
x_PM_NOR4xp25_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NOR4xp25_ASAP7_75t_R%noxref_14
cc_14 N_noxref_14_1 N_MM0_g 0.00159972f
cc_15 N_noxref_14_1 N_Y_16 0.0379781f
cc_16 N_noxref_14_1 N_noxref_13_1 0.00189464f
x_PM_NOR4xp25_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NOR4xp25_ASAP7_75t_R%noxref_13
cc_17 N_noxref_13_1 N_MM0_g 0.00351366f
cc_18 N_noxref_13_1 N_Y_15 0.0286725f
x_PM_NOR4xp25_ASAP7_75t_R%D VSS D N_MM3_g N_D_1 N_D_4 PM_NOR4xp25_ASAP7_75t_R%D
x_PM_NOR4xp25_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 N_C_4 PM_NOR4xp25_ASAP7_75t_R%C
cc_19 N_C_1 N_D_1 0.00150061f
cc_20 N_C_4 N_D_4 0.00661377f
cc_21 N_MM2_g N_MM3_g 0.00856971f
x_PM_NOR4xp25_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4 PM_NOR4xp25_ASAP7_75t_R%B
cc_22 N_B_1 N_C_1 0.00148896f
cc_23 N_B_4 N_C_4 0.00645733f
cc_24 N_MM1_g N_MM2_g 0.00869632f
x_PM_NOR4xp25_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM2_d N_MM1_d N_MM0_d N_MM7_d N_Y_1
+ N_Y_17 N_Y_13 N_Y_2 N_Y_14 N_Y_4 N_Y_19 N_Y_3 N_Y_16 N_Y_15 N_Y_18
+ PM_NOR4xp25_ASAP7_75t_R%Y
cc_25 N_Y_1 N_MM3_g 0.000860009f
cc_26 N_Y_17 N_D_4 0.00133602f
cc_27 N_Y_1 N_D_4 0.00192798f
cc_28 N_Y_13 N_MM3_g 0.0256833f
cc_29 N_Y_2 N_MM2_g 0.000716356f
cc_30 N_Y_17 N_C_4 0.00118791f
cc_31 N_Y_2 N_C_4 0.00175312f
cc_32 N_Y_14 N_MM2_g 0.0255737f
cc_33 N_Y_4 N_MM1_g 0.000355113f
cc_34 N_Y_2 N_MM1_g 0.000706172f
cc_35 N_Y_17 N_B_4 0.0011608f
cc_36 N_Y_4 N_B_4 0.00208553f
cc_37 N_Y_14 N_MM1_g 0.0265076f
cc_38 N_Y_19 N_A_4 0.000525554f
cc_39 N_Y_4 N_A_1 0.00073687f
cc_40 N_Y_3 N_MM0_g 0.000768811f
cc_41 N_Y_17 N_A_4 0.00111794f
cc_42 N_Y_16 N_A_1 0.00120666f
cc_43 N_Y_4 N_MM0_g 0.00169557f
cc_44 N_Y_15 N_MM0_g 0.010783f
cc_45 N_Y_18 N_A_4 0.00808823f
cc_46 N_Y_16 N_MM0_g 0.0498581f
*END of NOR4xp25_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR4xp75_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR4xp75_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR4xp75_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR4xp75_ASAP7_75t_R%PD2 VSS 16 17 29 30 33 34 10 13 1 11 12 3 2
c1 1 VSS 0.0030044f
c2 2 VSS 0.00310533f
c3 3 VSS 0.00301702f
c4 10 VSS 0.00209335f
c5 11 VSS 0.00206821f
c6 12 VSS 0.0020439f
c7 13 VSS 0.00316379f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 3 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r6 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r8 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r9 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4850 $Y2=0.1980
r10 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r11 24 25 9.56078 $w=1.3e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4440
+ $Y=0.1980 $X2=0.4850 $Y2=0.1980
r12 23 24 10.3769 $w=1.3e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3995
+ $Y=0.1980 $X2=0.4440 $Y2=0.1980
r13 22 23 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3995 $Y2=0.1980
r14 21 22 5.47996 $w=1.3e-08 $l=2.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3545
+ $Y=0.1980 $X2=0.3780 $Y2=0.1980
r15 20 21 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3230
+ $Y=0.1980 $X2=0.3545 $Y2=0.1980
r16 19 20 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2925
+ $Y=0.1980 $X2=0.3230 $Y2=0.1980
r17 18 19 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2925 $Y2=0.1980
r18 13 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1980 $X2=0.2700 $Y2=0.1980
r19 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r22 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r23 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0322822f
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0420294f
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%PD3 VSS 16 17 28 29 32 33 10 1 11 12 3 13 2
c1 1 VSS 0.0101252f
c2 2 VSS 0.00732232f
c3 3 VSS 0.00458479f
c4 10 VSS 0.00454341f
c5 11 VSS 0.00329097f
c6 12 VSS 0.00213718f
c7 13 VSS 0.0227404f
r1 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r2 3 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r4 32 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r5 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r6 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r8 28 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r9 3 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r10 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r11 23 24 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r12 22 23 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2405
+ $Y=0.2340 $X2=0.2855 $Y2=0.2340
r13 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2405 $Y2=0.2340
r14 20 21 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r15 19 20 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r16 18 19 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r17 13 18 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0935
+ $Y=0.2340 $X2=0.0970 $Y2=0.2340
r18 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r21 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r22 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0316126f
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00571356f
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%C VSS 7 3 4 5 8 1 6 9
c1 1 VSS 0.0119455f
c2 3 VSS 0.0367235f
c3 4 VSS 0.0368131f
c4 5 VSS 0.036851f
c5 6 VSS 0.0054214f
c6 7 VSS 0.00656004f
c7 8 VSS 0.0059828f
c8 9 VSS 0.00497072f
r1 8 28 4.53284 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.1600 $X2=0.2405 $Y2=0.1600
r2 6 9 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1600 $X2=0.2970 $Y2=0.1600
r3 6 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2720
+ $Y=0.1600 $X2=0.2405 $Y2=0.1600
r4 9 26 1.26576 $w=2.0056e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1600 $X2=0.2970 $Y2=0.1475
r5 5 22 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 7 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r7 7 26 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1475
r8 4 16 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 20 22 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r10 19 20 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r11 17 19 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r12 16 17 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r13 14 16 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r14 13 14 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r15 12 13 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r16 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r17 1 11 4.63801 $w=1.7681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r18 1 12 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r19 3 11 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r20 3 12 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%A VSS 20 3 4 5 1 6
c1 1 VSS 0.0151483f
c2 3 VSS 0.0383041f
c3 4 VSS 0.0382975f
c4 5 VSS 0.0383813f
c5 6 VSS 0.00817713f
r1 5 18 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r2 3 12 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 20 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.0980
r4 16 18 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r5 15 16 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r6 14 15 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r7 10 12 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5795 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r8 9 10 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.5940
+ $Y=0.1350 $X2=0.5795 $Y2=0.1350
r9 8 9 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.6085
+ $Y=0.1350 $X2=0.5940 $Y2=0.1350
r10 4 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r11 20 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
r12 4 8 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6085 $Y2=0.1350
r13 4 14 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%PD1 VSS 16 17 29 30 33 34 10 1 13 11 3 12 2
c1 1 VSS 0.0047093f
c2 2 VSS 0.00418584f
c3 3 VSS 0.00449435f
c4 10 VSS 0.0021652f
c5 11 VSS 0.00208567f
c6 12 VSS 0.00214859f
c7 13 VSS 0.0217837f
r1 34 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r2 3 32 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6480 $Y2=0.2025
r4 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r5 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r6 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r7 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r8 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r9 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.2340
r10 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r11 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6095
+ $Y=0.2340 $X2=0.6480 $Y2=0.2340
r12 23 24 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5645
+ $Y=0.2340 $X2=0.6095 $Y2=0.2340
r13 22 23 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5645 $Y2=0.2340
r14 21 22 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5175
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r15 20 21 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.5015
+ $Y=0.2340 $X2=0.5175 $Y2=0.2340
r16 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4700
+ $Y=0.2340 $X2=0.5015 $Y2=0.2340
r17 18 19 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4700 $Y2=0.2340
r18 13 18 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.4175
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r19 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r22 10 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r23 16 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%D VSS 28 3 4 5 1 11 8 9
c1 1 VSS 0.00936162f
c2 3 VSS 0.0704347f
c3 4 VSS 0.0700172f
c4 5 VSS 0.0697732f
c5 6 VSS 0.0121676f
c6 7 VSS 0.0118696f
c7 8 VSS 0.00508181f
c8 9 VSS 0.0103502f
c9 10 VSS 0.00322911f
c10 11 VSS 0.0102691f
r1 11 38 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r2 9 35 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r3 37 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2035 $X2=0.0270 $Y2=0.2160
r4 36 37 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1755 $X2=0.0270 $Y2=0.2035
r5 7 10 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1475 $X2=0.0270 $Y2=0.1350
r6 7 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1475 $X2=0.0270 $Y2=0.1755
r7 6 10 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0980 $X2=0.0270 $Y2=0.1350
r8 6 35 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0980 $X2=0.0270 $Y2=0.0575
r9 10 30 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1350 $X2=0.0465 $Y2=0.1350
r10 5 26 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r11 4 20 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r12 28 8 3.84763 $w=1.3e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0645 $Y2=0.1350
r13 8 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0645
+ $Y=0.1350 $X2=0.0465 $Y2=0.1350
r14 24 26 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r15 23 24 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r16 21 23 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r17 20 21 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r18 18 20 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r19 17 18 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r20 16 17 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r21 14 16 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r22 13 14 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r23 28 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r24 1 13 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r25 1 15 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r26 3 13 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r27 3 15 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r28 3 16 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%B VSS 27 3 4 5 8 7 1 6
c1 1 VSS 0.0133591f
c2 3 VSS 0.0374375f
c3 4 VSS 0.0373138f
c4 5 VSS 0.0372942f
c5 6 VSS 0.00704992f
c6 7 VSS 0.005572f
c7 8 VSS 0.0059744f
r1 8 30 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.1575 $X2=0.5400 $Y2=0.1665
r2 29 30 1.30447 $w=1.47857e-08 $l=1.49833e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5265 $Y=0.1600 $X2=0.5400 $Y2=0.1665
r3 7 28 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1600 $X2=0.5130 $Y2=0.1475
r4 7 29 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1600 $X2=0.5265 $Y2=0.1600
r5 27 28 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1475
r6 27 6 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.0980
r7 5 22 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r8 4 15 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r9 27 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r10 21 22 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r11 19 21 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5035 $Y2=0.1350
r12 18 19 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r13 16 18 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r14 15 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r15 13 15 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r16 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r17 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r18 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r19 1 10 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r20 1 11 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r21 3 10 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r22 3 11 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_NOR4xp75_ASAP7_75t_R%Y VSS 80 40 41 65 66 69 70 73 74 77 78 85 86 95
+ 98 99 33 26 1 2 25 3 27 5 29 4 28 34 32 6 30 8 35 7 31
c1 1 VSS 0.00877771f
c2 2 VSS 0.00878609f
c3 3 VSS 0.00872445f
c4 4 VSS 0.00848472f
c5 5 VSS 0.00814813f
c6 6 VSS 0.00280616f
c7 7 VSS 0.00814167f
c8 8 VSS 0.00414188f
c9 25 VSS 0.00396939f
c10 26 VSS 0.00391197f
c11 27 VSS 0.00389571f
c12 28 VSS 0.00385302f
c13 29 VSS 0.00384858f
c14 30 VSS 0.00379713f
c15 31 VSS 0.00210266f
c16 32 VSS 0.0023091f
c17 33 VSS 0.0571292f
c18 34 VSS 0.00175749f
c19 35 VSS 0.00374907f
c20 36 VSS 0.00338938f
c21 37 VSS 0.00105773f
r1 99 97 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r2 6 97 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r3 31 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5940 $Y2=0.2025
r4 98 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r5 32 8 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.2025 $X2=0.7000 $Y2=0.2025
r6 95 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.2025 $X2=0.6875 $Y2=0.2025
r7 6 92 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.1980
r8 8 87 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.2025
+ $X2=0.7030 $Y2=0.1980
r9 92 93 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.1980 $X2=0.6075 $Y2=0.1980
r10 90 93 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1980 $X2=0.6075 $Y2=0.1980
r11 89 90 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.1980 $X2=0.6210 $Y2=0.1980
r12 87 88 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.7030
+ $Y=0.1980 $X2=0.7160 $Y2=0.1980
r13 34 87 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.6800
+ $Y=0.1980 $X2=0.7030 $Y2=0.1980
r14 34 89 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6800
+ $Y=0.1980 $X2=0.6480 $Y2=0.1980
r15 37 82 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1765
r16 37 88 1.38235 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7160 $Y2=0.1980
r17 86 84 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0540 $X2=0.6625 $Y2=0.0540
r18 7 84 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.0540 $X2=0.6625 $Y2=0.0540
r19 30 7 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0540 $X2=0.6480 $Y2=0.0540
r20 85 30 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0540 $X2=0.6335 $Y2=0.0540
r21 81 82 4.95528 $w=1.3e-08 $l=2.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1552 $X2=0.7290 $Y2=0.1765
r22 80 81 2.15701 $w=1.3e-08 $l=9.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1460 $X2=0.7290 $Y2=0.1552
r23 80 79 8.91951 $w=1.3e-08 $l=3.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1460 $X2=0.7290 $Y2=0.1077
r24 35 36 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0575 $X2=0.7290 $Y2=0.0360
r25 35 79 11.7178 $w=1.3e-08 $l=5.02e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.0575 $X2=0.7290 $Y2=0.1077
r26 78 76 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0540 $X2=0.5545 $Y2=0.0540
r27 5 76 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0540 $X2=0.5545 $Y2=0.0540
r28 29 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0540 $X2=0.5400 $Y2=0.0540
r29 77 29 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0540 $X2=0.5255 $Y2=0.0540
r30 74 72 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0540 $X2=0.4465 $Y2=0.0540
r31 4 72 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0540 $X2=0.4465 $Y2=0.0540
r32 28 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0540 $X2=0.4320 $Y2=0.0540
r33 73 28 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0540 $X2=0.4175 $Y2=0.0540
r34 70 68 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0540 $X2=0.3385 $Y2=0.0540
r35 3 68 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0540 $X2=0.3385 $Y2=0.0540
r36 27 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3240 $Y2=0.0540
r37 69 27 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r38 66 64 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r39 2 64 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r40 26 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r41 65 26 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r42 7 61 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0540
+ $X2=0.6480 $Y2=0.0360
r43 36 62 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.0360 $X2=0.6885 $Y2=0.0360
r44 5 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0540
+ $X2=0.5400 $Y2=0.0360
r45 4 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0540
+ $X2=0.4320 $Y2=0.0360
r46 3 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r47 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r48 61 62 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6885 $Y2=0.0360
r49 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r50 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6345 $Y2=0.0360
r51 58 59 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5960
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r52 57 58 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5645
+ $Y=0.0360 $X2=0.5960 $Y2=0.0360
r53 56 57 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5645 $Y2=0.0360
r54 55 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r55 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5265 $Y2=0.0360
r56 53 54 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5015
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r57 52 53 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4700
+ $Y=0.0360 $X2=0.5015 $Y2=0.0360
r58 51 52 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4700 $Y2=0.0360
r59 50 51 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r60 49 50 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r61 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r62 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r63 46 47 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r64 45 46 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r65 44 45 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r66 43 44 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r67 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r68 33 42 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.0970 $Y2=0.0360
r69 1 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r70 41 39 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r71 1 39 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r72 25 1 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r73 40 25 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
.ends


*
.SUBCKT NOR4xp75_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3@3 N_MM3@3_d N_MM4@3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3@2 N_MM3@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2@3 N_MM2@3_d N_MM5@3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2@2 N_MM2@2_d N_MM5@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@3 N_MM1@3_d N_MM6@3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 N_MM1@2_d N_MM6@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@3 N_MM0@3_d N_MM0@3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM4@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 N_MM5@3_d N_MM5@3_g N_MM5@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM5@2_g N_MM5@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@3 N_MM6@3_d N_MM6@3_g N_MM6@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g N_MM6@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@3 N_MM7@3_d N_MM0@3_g N_MM7@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM0@2_g N_MM7@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR4xp75_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR4xp75_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR4xp75_ASAP7_75t_R%PD2 VSS N_MM5_d N_MM5@3_d N_MM5@2_d N_MM6_s N_MM6@3_s
+ N_MM6@2_s N_PD2_10 N_PD2_13 N_PD2_1 N_PD2_11 N_PD2_12 N_PD2_3 N_PD2_2
+ PM_NOR4xp75_ASAP7_75t_R%PD2
cc_1 N_PD2_10 N_C_8 0.000484268f
cc_2 N_PD2_10 N_MM5@2_g 0.000726601f
cc_3 N_PD2_13 N_C_6 0.00166528f
cc_4 N_PD2_1 N_MM5_g 0.00187353f
cc_5 N_PD2_10 N_C_1 0.00290973f
cc_6 N_PD2_13 N_C_9 0.00408076f
cc_7 N_PD2_11 N_MM5@2_g 0.0325029f
cc_8 N_PD2_10 N_MM5@3_g 0.0180004f
cc_9 N_PD2_10 N_MM5_g 0.0491199f
cc_10 N_PD2_12 N_MM6_g 0.000739626f
cc_11 N_PD2_12 N_B_7 0.000776821f
cc_12 N_PD2_13 N_B_1 0.00154714f
cc_13 N_PD2_3 N_MM6@3_g 0.00179719f
cc_14 N_PD2_12 N_B_1 0.00363567f
cc_15 N_PD2_11 N_MM6_g 0.0325291f
cc_16 N_PD2_12 N_MM6@2_g 0.0179411f
cc_17 N_PD2_12 N_MM6@3_g 0.049757f
cc_18 N_PD2_10 N_PD3_13 0.00110095f
cc_19 N_PD2_10 N_PD3_11 0.00110424f
cc_20 N_PD2_2 N_PD3_3 0.00126019f
cc_21 N_PD2_1 N_PD3_3 0.00301873f
cc_22 N_PD2_1 N_PD3_2 0.00399228f
cc_23 N_PD2_13 N_PD3_13 0.0116845f
x_PM_NOR4xp75_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_NOR4xp75_ASAP7_75t_R%noxref_11
cc_24 N_noxref_11_1 N_MM3_g 0.00448205f
x_PM_NOR4xp75_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_NOR4xp75_ASAP7_75t_R%noxref_12
cc_25 N_noxref_12_1 N_MM3_g 0.00247244f
cc_26 N_noxref_12_1 N_noxref_11_1 0.00189547f
x_PM_NOR4xp75_ASAP7_75t_R%PD3 VSS N_MM4_d N_MM4@3_d N_MM4@2_d N_MM5_s N_MM5@3_s
+ N_MM5@2_s N_PD3_10 N_PD3_1 N_PD3_11 N_PD3_12 N_PD3_3 N_PD3_13 N_PD3_2
+ PM_NOR4xp75_ASAP7_75t_R%PD3
cc_27 N_PD3_10 N_MM4@2_g 0.00208831f
cc_28 N_PD3_10 N_D_11 0.000460652f
cc_29 N_PD3_1 N_MM3_g 0.00195342f
cc_30 N_PD3_10 N_D_1 0.0028693f
cc_31 N_PD3_11 N_MM4@2_g 0.0328386f
cc_32 N_PD3_10 N_MM4@3_g 0.0181767f
cc_33 N_PD3_10 N_MM3_g 0.0494159f
cc_34 N_PD3_12 N_MM5_g 0.00183683f
cc_35 N_PD3_3 N_MM5@3_g 0.00184703f
cc_36 N_PD3_12 N_C_1 0.00259096f
cc_37 N_PD3_13 N_C_8 0.00308097f
cc_38 N_PD3_11 N_MM5_g 0.0328671f
cc_39 N_PD3_12 N_MM5@2_g 0.0180983f
cc_40 N_PD3_12 N_MM5@3_g 0.0496053f
x_PM_NOR4xp75_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NOR4xp75_ASAP7_75t_R%noxref_13
cc_41 N_noxref_13_1 N_MM0@2_g 0.00348273f
cc_42 N_noxref_13_1 N_Y_35 0.000356772f
cc_43 N_noxref_13_1 N_Y_30 0.00123434f
x_PM_NOR4xp75_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NOR4xp75_ASAP7_75t_R%noxref_14
cc_44 N_noxref_14_1 N_MM0@2_g 0.00160127f
cc_45 N_noxref_14_1 N_Y_8 0.00049461f
cc_46 N_noxref_14_1 N_Y_32 0.0366785f
cc_47 N_noxref_14_1 N_noxref_13_1 0.00188936f
x_PM_NOR4xp75_ASAP7_75t_R%C VSS C N_MM5_g N_MM5@3_g N_MM5@2_g N_C_8 N_C_1 N_C_6
+ N_C_9 PM_NOR4xp75_ASAP7_75t_R%C
cc_48 N_C_8 N_D_1 0.00148265f
cc_49 N_MM5_g N_MM4@2_g 0.00675473f
x_PM_NOR4xp75_ASAP7_75t_R%A VSS A N_MM7_g N_MM0@3_g N_MM0@2_g N_A_1 N_A_6
+ PM_NOR4xp75_ASAP7_75t_R%A
cc_50 N_A_1 N_B_8 0.00159343f
cc_51 N_MM7_g N_MM6@2_g 0.00753392f
x_PM_NOR4xp75_ASAP7_75t_R%PD1 VSS N_MM6_d N_MM6@3_d N_MM6@2_d N_MM7_s N_MM7@3_s
+ N_MM7@2_s N_PD1_10 N_PD1_1 N_PD1_13 N_PD1_11 N_PD1_3 N_PD1_12 N_PD1_2
+ PM_NOR4xp75_ASAP7_75t_R%PD1
cc_52 N_PD1_10 N_MM6@2_g 0.0014133f
cc_53 N_PD1_1 N_MM6_g 0.00172315f
cc_54 N_PD1_13 N_B_8 0.00249f
cc_55 N_PD1_10 N_B_1 0.00304711f
cc_56 N_PD1_11 N_MM6@2_g 0.0329886f
cc_57 N_PD1_10 N_MM6@3_g 0.0182386f
cc_58 N_PD1_10 N_MM6_g 0.0499434f
cc_59 N_PD1_3 N_MM0@3_g 0.0017623f
cc_60 N_PD1_12 N_A_1 0.00276462f
cc_61 N_PD1_11 N_MM7_g 0.0329709f
cc_62 N_PD1_12 N_MM0@2_g 0.0181927f
cc_63 N_PD1_12 N_MM0@3_g 0.0500592f
cc_64 N_PD1_10 N_PD2_11 0.00110359f
cc_65 N_PD1_10 N_PD2_12 0.00110472f
cc_66 N_PD1_2 N_PD2_3 0.00125863f
cc_67 N_PD1_1 N_PD2_3 0.00273371f
cc_68 N_PD1_1 N_PD2_2 0.00443369f
cc_69 N_PD1_13 N_PD2_13 0.0121872f
x_PM_NOR4xp75_ASAP7_75t_R%D VSS D N_MM3_g N_MM4@3_g N_MM4@2_g N_D_1 N_D_11
+ N_D_8 N_D_9 PM_NOR4xp75_ASAP7_75t_R%D
x_PM_NOR4xp75_ASAP7_75t_R%B VSS B N_MM6_g N_MM6@3_g N_MM6@2_g N_B_8 N_B_7 N_B_1
+ N_B_6 PM_NOR4xp75_ASAP7_75t_R%B
cc_70 N_MM6_g N_MM5@2_g 0.00710587f
x_PM_NOR4xp75_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM3@3_d N_MM3@2_d N_MM2_d N_MM2@3_d
+ N_MM2@2_d N_MM1_d N_MM1@3_d N_MM1@2_d N_MM0_d N_MM0@3_d N_MM0@2_d N_MM7@2_d
+ N_MM7_d N_MM7@3_d N_Y_33 N_Y_26 N_Y_1 N_Y_2 N_Y_25 N_Y_3 N_Y_27 N_Y_5 N_Y_29
+ N_Y_4 N_Y_28 N_Y_34 N_Y_32 N_Y_6 N_Y_30 N_Y_8 N_Y_35 N_Y_7 N_Y_31
+ PM_NOR4xp75_ASAP7_75t_R%Y
cc_71 N_Y_33 N_MM3_g 0.000334349f
cc_72 N_Y_26 N_MM3_g 0.000349758f
cc_73 N_Y_1 N_D_8 0.000380944f
cc_74 N_Y_33 N_D_9 0.000440358f
cc_75 N_Y_2 N_MM4@2_g 0.00052479f
cc_76 N_Y_33 N_MM4@2_g 0.00109039f
cc_77 N_Y_1 N_MM3_g 0.00117557f
cc_78 N_Y_25 N_D_1 0.0011829f
cc_79 N_Y_26 N_MM4@2_g 0.0240417f
cc_80 N_Y_25 N_MM4@3_g 0.0134135f
cc_81 N_Y_25 N_MM3_g 0.0360312f
cc_82 N_Y_3 N_MM5@3_g 0.0013559f
cc_83 N_Y_2 N_MM5@3_g 0.000490744f
cc_84 N_Y_26 N_MM5@3_g 0.000331716f
cc_85 N_Y_2 N_MM5_g 0.000591718f
cc_86 N_Y_27 N_C_1 0.00107477f
cc_87 N_Y_3 N_C 0.00213009f
cc_88 N_Y_33 N_C 0.00215917f
cc_89 N_Y_26 N_MM5_g 0.0239925f
cc_90 N_Y_27 N_MM5@2_g 0.0133893f
cc_91 N_Y_27 N_MM5@3_g 0.035939f
cc_92 N_Y_5 N_MM6_g 0.000375991f
cc_93 N_Y_33 N_MM6_g 0.00018289f
cc_94 N_Y_29 N_MM6_g 0.000349762f
cc_95 N_Y_5 N_MM6@2_g 0.000755644f
cc_96 N_Y_4 N_MM6_g 0.00100921f
cc_97 N_Y_28 N_B_1 0.00125465f
cc_98 N_Y_34 N_B_8 0.00151643f
cc_99 N_Y_33 N_B_6 0.00179904f
cc_100 N_Y_5 N_B_6 0.00226637f
cc_101 N_Y_29 N_MM6@2_g 0.0241282f
cc_102 N_Y_28 N_MM6@3_g 0.0134365f
cc_103 N_Y_28 N_MM6_g 0.0359745f
cc_104 N_Y_29 N_MM7_g 0.0109216f
cc_105 N_Y_32 N_MM7_g 0.000471513f
cc_106 N_Y_6 N_MM7_g 0.00232741f
cc_107 N_Y_5 N_MM7_g 0.000530761f
cc_108 N_Y_30 N_MM0@3_g 0.0220575f
cc_109 N_Y_8 N_MM0@2_g 0.000854822f
cc_110 N_Y_35 N_A_1 0.000903187f
cc_111 N_Y_7 N_MM0@3_g 0.00126458f
cc_112 N_Y_34 N_A_6 0.00163547f
cc_113 N_Y_33 N_A_6 0.00168463f
cc_114 N_Y_7 N_A_6 0.00401318f
cc_115 N_Y_31 N_A_1 0.00470215f
cc_116 N_Y_32 N_MM0@2_g 0.0471025f
cc_117 N_Y_31 N_MM0@3_g 0.0319106f
cc_118 N_Y_31 N_MM7_g 0.0633607f
cc_119 N_Y_6 N_PD1_13 0.000831688f
cc_120 N_Y_8 N_PD1_13 0.000242346f
cc_121 N_Y_32 N_PD1_13 0.000555487f
cc_122 N_Y_31 N_PD1_13 0.000567824f
cc_123 N_Y_31 N_PD1_11 0.00110975f
cc_124 N_Y_31 N_PD1_12 0.00112749f
cc_125 N_Y_8 N_PD1_3 0.00128985f
cc_126 N_Y_6 N_PD1_3 0.00316918f
cc_127 N_Y_6 N_PD1_2 0.00408636f
cc_128 N_Y_34 N_PD1_13 0.0101049f
*END of NOR4xp75_ASAP7_75t_R.pxi
.ENDS
** Design:	NOR5xp2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "NOR5xp2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "NOR5xp2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_NOR5xp2_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000849971f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0425574f
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000889469f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%NET024 VSS 2 3 1
c1 1 VSS 0.000879335f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%NET023 VSS 2 3 1
c1 1 VSS 0.00084846f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%E VSS 8 3 1 4
c1 1 VSS 0.00365915f
c2 3 VSS 0.0714757f
c3 4 VSS 0.0151516f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1360 $X2=0.2970 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1360
+ $X2=0.2970 $Y2=0.1355
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00550086f
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%D VSS 8 3 1 4
c1 1 VSS 0.00405293f
c2 3 VSS 0.0354821f
c3 4 VSS 0.00718881f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1360 $X2=0.2430 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1360
+ $X2=0.2430 $Y2=0.1355
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00401944f
c2 3 VSS 0.0351111f
c3 4 VSS 0.00688582f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1360
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00418386f
c2 3 VSS 0.0353074f
c3 4 VSS 0.00729743f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1360 $X2=0.1890 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1360
+ $X2=0.1890 $Y2=0.1355
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0316565f
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00513957f
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%A VSS 11 3 1 4
c1 1 VSS 0.0055569f
c2 3 VSS 0.0349871f
c3 4 VSS 0.00434373f
r1 11 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0810 $Y2=0.0985
r2 7 10 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1360 $X2=0.0915 $Y2=0.1360
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0905 $Y2=0.1360
r4 11 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1360
+ $X2=0.0810 $Y2=0.1360
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0810 $Y2=0.1360
r6 1 8 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0685 $Y2=0.1360
r7 3 6 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1360
r8 3 8 4.17867 $w=1.8386e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1360
r9 3 10 1.08747 $w=2.16729e-07 $l=1.05475e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1360
.ends

.subckt PM_NOR5xp2_ASAP7_75t_R%Y VSS 43 23 24 48 49 51 56 20 2 1 18 16 13 17 3
+ 14 4 15
c1 1 VSS 0.0060518f
c2 2 VSS 0.0085602f
c3 3 VSS 0.00845254f
c4 4 VSS 0.00751471f
c5 13 VSS 0.00388946f
c6 14 VSS 0.00389842f
c7 15 VSS 0.00337714f
c8 16 VSS 0.00261731f
c9 17 VSS 0.0042531f
c10 18 VSS 0.0292837f
c11 19 VSS 0.00333914f
c12 20 VSS 0.00601286f
r1 56 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 16 55 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 1 53 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 52 53 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0410
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 20 45 3.31868 $w=1.62766e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2115
r6 20 52 1.9532 $w=1.65714e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0410 $Y2=0.2340
r7 15 4 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0540 $X2=0.3220 $Y2=0.0540
r8 51 15 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0540 $X2=0.3095 $Y2=0.0540
r9 49 47 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r10 3 47 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r11 14 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r12 48 14 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r13 44 45 7.10752 $w=1.5e-08 $l=4.18e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1697 $X2=0.0270 $Y2=0.2115
r14 43 44 4.8944 $w=1.5e-08 $l=2.87e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1410 $X2=0.0270 $Y2=0.1697
r15 43 42 6.08608 $w=1.5e-08 $l=3.58e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1410 $X2=0.0270 $Y2=0.1052
r16 17 19 2.56637 $w=1.7093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r17 17 42 8.12896 $w=1.5e-08 $l=4.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1052
r18 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0540
+ $X2=0.3240 $Y2=0.0360
r19 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r20 19 29 4.28601 $w=1.71509e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0535 $Y2=0.0360
r21 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r22 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r23 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r24 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r25 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r26 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r27 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r28 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r29 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 30 31 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r31 28 29 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0710
+ $Y=0.0360 $X2=0.0535 $Y2=0.0360
r32 27 28 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0710 $Y2=0.0360
r33 26 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r34 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r35 18 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r36 18 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r37 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r38 24 22 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r39 2 22 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r40 13 2 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r41 23 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r42 1 16 1e-05
.ends


*
.SUBCKT NOR5xp2_ASAP7_75t_R VSS VDD A B C D E Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* E E
* Y Y
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM0_g N_MM9_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM1_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM2_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM3_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "NOR5xp2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "NOR5xp2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_NOR5xp2_ASAP7_75t_R%NET30 VSS N_MM7_s N_MM6_d N_NET30_1
+ PM_NOR5xp2_ASAP7_75t_R%NET30
cc_1 N_NET30_1 N_MM2_g 0.0174606f
cc_2 N_NET30_1 N_MM3_g 0.0175648f
x_PM_NOR5xp2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_NOR5xp2_ASAP7_75t_R%noxref_16
cc_3 N_noxref_16_1 N_MM4_g 0.00185555f
cc_4 N_noxref_16_1 N_noxref_15_1 0.00192724f
x_PM_NOR5xp2_ASAP7_75t_R%NET29 VSS N_MM6_s N_MM5_d N_NET29_1
+ PM_NOR5xp2_ASAP7_75t_R%NET29
cc_5 N_NET29_1 N_MM3_g 0.0172585f
cc_6 N_NET29_1 N_MM4_g 0.0172476f
x_PM_NOR5xp2_ASAP7_75t_R%NET024 VSS N_MM9_s N_MM8_d N_NET024_1
+ PM_NOR5xp2_ASAP7_75t_R%NET024
cc_7 N_NET024_1 N_MM0_g 0.0172318f
cc_8 N_NET024_1 N_MM1_g 0.0172857f
x_PM_NOR5xp2_ASAP7_75t_R%NET023 VSS N_MM8_s N_MM7_d N_NET023_1
+ PM_NOR5xp2_ASAP7_75t_R%NET023
cc_9 N_NET023_1 N_MM1_g 0.0174588f
cc_10 N_NET023_1 N_MM2_g 0.017568f
x_PM_NOR5xp2_ASAP7_75t_R%E VSS E N_MM4_g N_E_1 N_E_4 PM_NOR5xp2_ASAP7_75t_R%E
cc_11 N_E_1 N_D_1 0.00164559f
cc_12 N_E_4 N_D_4 0.0068765f
cc_13 N_MM4_g N_MM3_g 0.00852147f
x_PM_NOR5xp2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_NOR5xp2_ASAP7_75t_R%noxref_15
cc_14 N_noxref_15_1 N_MM4_g 0.00374019f
cc_15 N_noxref_15_1 N_Y_15 0.0273439f
x_PM_NOR5xp2_ASAP7_75t_R%D VSS D N_MM3_g N_D_1 N_D_4 PM_NOR5xp2_ASAP7_75t_R%D
cc_16 N_D_1 N_C_1 0.00169547f
cc_17 N_D_4 N_C_4 0.00637701f
cc_18 N_MM3_g N_MM2_g 0.00866575f
x_PM_NOR5xp2_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4 PM_NOR5xp2_ASAP7_75t_R%B
cc_19 N_B_1 N_A_1 0.00152283f
cc_20 N_B_4 N_A_4 0.00525842f
cc_21 N_MM1_g N_MM0_g 0.00837488f
x_PM_NOR5xp2_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 N_C_4 PM_NOR5xp2_ASAP7_75t_R%C
cc_22 N_C_1 N_B_1 0.00165584f
cc_23 N_C_4 N_B_4 0.00642113f
cc_24 N_MM2_g N_MM1_g 0.00869612f
x_PM_NOR5xp2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_NOR5xp2_ASAP7_75t_R%noxref_13
cc_25 N_noxref_13_1 N_MM0_g 0.00358771f
cc_26 N_noxref_13_1 N_Y_13 0.00151893f
x_PM_NOR5xp2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_NOR5xp2_ASAP7_75t_R%noxref_14
cc_27 N_noxref_14_1 N_MM0_g 0.00166236f
cc_28 N_noxref_14_1 N_Y_16 0.037818f
cc_29 N_noxref_14_1 N_noxref_13_1 0.0018885f
x_PM_NOR5xp2_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_NOR5xp2_ASAP7_75t_R%A
x_PM_NOR5xp2_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM1_d N_MM2_d N_MM3_d N_MM4_d
+ N_MM9_d N_Y_20 N_Y_2 N_Y_1 N_Y_18 N_Y_16 N_Y_13 N_Y_17 N_Y_3 N_Y_14 N_Y_4
+ N_Y_15 PM_NOR5xp2_ASAP7_75t_R%Y
cc_30 N_Y_20 N_A_4 0.000512512f
cc_31 N_Y_2 N_MM0_g 0.000662139f
cc_32 N_Y_1 N_A_1 0.000686532f
cc_33 N_Y_18 N_A_4 0.00110305f
cc_34 N_Y_16 N_A_1 0.00168509f
cc_35 N_Y_1 N_MM0_g 0.00193005f
cc_36 N_Y_13 N_MM0_g 0.0108466f
cc_37 N_Y_17 N_A_4 0.00812079f
cc_38 N_Y_16 N_MM0_g 0.0497476f
cc_39 N_Y_1 N_MM1_g 0.000346001f
cc_40 N_Y_2 N_MM1_g 0.000701136f
cc_41 N_Y_18 N_B_4 0.00118412f
cc_42 N_Y_1 N_B_4 0.002101f
cc_43 N_Y_13 N_MM1_g 0.0265138f
cc_44 N_Y_3 N_MM2_g 0.000672299f
cc_45 N_Y_18 N_C_4 0.00122001f
cc_46 N_Y_3 N_C_4 0.00160187f
cc_47 N_Y_14 N_MM2_g 0.0254933f
cc_48 N_Y_3 N_MM3_g 0.00066683f
cc_49 N_Y_18 N_D_4 0.00123607f
cc_50 N_Y_3 N_D_4 0.00166773f
cc_51 N_Y_14 N_MM3_g 0.0254751f
cc_52 N_Y_4 N_MM4_g 0.000851013f
cc_53 N_Y_18 N_E_4 0.00132528f
cc_54 N_Y_4 N_E_4 0.00187922f
cc_55 N_Y_15 N_MM4_g 0.0256037f
*END of NOR5xp2_ASAP7_75t_R.pxi
.ENDS
** Design:	AND2x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND2x2_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00497172f
.ends

.subckt PM_AND2x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0422936f
.ends

.subckt PM_AND2x2_ASAP7_75t_R%A VSS 4 3 1
c1 1 VSS 0.0055481f
c2 3 VSS 0.0825682f
c3 4 VSS 0.00381638f
r1 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AND2x2_ASAP7_75t_R%NET20 VSS 2 3 1
c1 1 VSS 0.000681943f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND2x2_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.031612f
.ends

.subckt PM_AND2x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0422379f
.ends

.subckt PM_AND2x2_ASAP7_75t_R%Y VSS 27 20 21 34 35 7 10 8 15 14 2 1 9
c1 1 VSS 0.00835707f
c2 2 VSS 0.00840842f
c3 7 VSS 0.00458009f
c4 8 VSS 0.00451005f
c5 9 VSS 0.00108144f
c6 10 VSS 0.00124187f
c7 11 VSS 0.00658603f
c8 12 VSS 0.00656171f
c9 13 VSS 0.00719591f
c10 14 VSS 0.00209353f
c11 15 VSS 0.00218018f
c12 16 VSS 0.00347703f
c13 17 VSS 0.00352861f
r1 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 2 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 34 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 2 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2160 $Y2=0.2160
r7 10 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1865 $X2=0.2160 $Y2=0.1980
r8 15 31 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2160 $Y2=0.2160
r9 12 17 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2565 $Y=0.2340 $X2=0.2970 $Y2=0.2340
r10 12 15 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2565 $Y=0.2340 $X2=0.2160 $Y2=0.2340
r11 17 29 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2970 $Y2=0.2045
r12 28 29 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1660 $X2=0.2970 $Y2=0.2045
r13 27 28 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1660
r14 27 26 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1455
r15 25 26 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1455
r16 24 25 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1060 $X2=0.2970 $Y2=0.1350
r17 13 16 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0655 $X2=0.2970 $Y2=0.0360
r18 13 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0655 $X2=0.2970 $Y2=0.1060
r19 11 14 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2565 $Y=0.0360 $X2=0.2160 $Y2=0.0360
r20 11 16 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2565 $Y=0.0360 $X2=0.2970 $Y2=0.0360
r21 9 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0720
r22 9 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0360
r23 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r24 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r25 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r26 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r27 20 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends

.subckt PM_AND2x2_ASAP7_75t_R%B VSS 14 3 1 6 4 5
c1 1 VSS 0.00146635f
c2 3 VSS 0.032528f
c3 4 VSS 0.00883551f
c4 5 VSS 0.0110316f
c5 6 VSS 0.00181483f
c6 7 VSS 0.00159436f
r1 5 7 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1720 $X2=0.0270 $Y2=0.1350
r2 4 7 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1060 $X2=0.0270 $Y2=0.1350
r3 14 6 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0655
+ $Y=0.1350 $X2=0.0485 $Y2=0.1350
r4 6 7 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0485
+ $Y=0.1350 $X2=0.0270 $Y2=0.1350
r5 1 9 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0750
+ $Y=0.1345 $X2=0.0850 $Y2=0.1345
r6 1 10 2.09261 $w=2.04231e-08 $l=6.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0750 $Y=0.1345 $X2=0.0685 $Y2=0.1345
r7 14 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0655 $Y=0.1350
+ $X2=0.0750 $Y2=0.1345
r8 3 9 1.73446 $w=1.505e-07 $l=4.03113e-09 $layer=LIG $thickness=5.3e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0850 $Y2=0.1345
r9 3 10 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1345
.ends

.subckt PM_AND2x2_ASAP7_75t_R%NET10 VSS 9 10 52 53 55 18 3 4 13 15 11 12 20 14
+ 1 17 16 21 19
c1 1 VSS 0.00797624f
c2 3 VSS 0.00806448f
c3 4 VSS 0.00913062f
c4 9 VSS 0.0803232f
c5 10 VSS 0.0808875f
c6 11 VSS 0.00678543f
c7 12 VSS 0.00748318f
c8 13 VSS 0.00165686f
c9 14 VSS 0.00855063f
c10 15 VSS 0.00860441f
c11 16 VSS 0.00315094f
c12 17 VSS 0.00316917f
c13 18 VSS 0.00317328f
c14 19 VSS 0.00301967f
c15 20 VSS 0.00103165f
c16 21 VSS 0.00299477f
r1 55 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r2 11 54 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r3 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0665 $Y=0.0675
+ $X2=0.0790 $Y2=0.0755
r4 53 51 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r5 4 51 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r6 12 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r7 52 12 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r8 47 48 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.0665 $X2=0.0790 $Y2=0.0755
r9 13 47 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.0540 $X2=0.0790 $Y2=0.0665
r10 13 46 2.65995 $w=1.48966e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0790 $Y=0.0540 $X2=0.0790 $Y2=0.0395
r11 4 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1080 $Y2=0.2340
r12 18 41 1.05672 $w=1.56923e-08 $l=1.32004e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0790 $Y=0.0305 $X2=0.0910 $Y2=0.0360
r13 18 46 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0790
+ $Y=0.0305 $X2=0.0790 $Y2=0.0395
r14 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r15 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r16 15 21 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1710 $Y2=0.2340
r17 15 42 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r18 40 41 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1100
+ $Y=0.0360 $X2=0.0910 $Y2=0.0360
r19 39 40 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1100 $Y2=0.0360
r20 14 19 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1710 $Y2=0.0360
r21 14 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r22 21 38 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.2340 $X2=0.1710 $Y2=0.2125
r23 19 36 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.0360 $X2=0.1710 $Y2=0.0575
r24 37 38 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1920 $X2=0.1710 $Y2=0.2125
r25 17 20 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.1640 $X2=0.1710 $Y2=0.1350
r26 17 37 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1640 $X2=0.1710 $Y2=0.1920
r27 35 36 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0780 $X2=0.1710 $Y2=0.0575
r28 16 20 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.1060 $X2=0.1710 $Y2=0.1350
r29 16 35 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1060 $X2=0.1710 $Y2=0.0780
r30 10 30 2.68099 $w=1.25e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1345
r31 20 32 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r32 28 30 3.5124 $w=2.166e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1345 $X2=0.2430 $Y2=0.1345
r33 27 28 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1345 $X2=0.2305 $Y2=0.1345
r34 26 27 6.64723 $w=1.63e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1345 $X2=0.2160 $Y2=0.1345
r35 24 26 1.26439 $w=1.74167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1985 $Y=0.1345 $X2=0.2015 $Y2=0.1345
r36 23 24 2.24801 $w=2.3e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1345 $X2=0.1985 $Y2=0.1345
r37 23 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1345
+ $X2=0.1890 $Y2=0.1350
r38 1 23 2.24801 $w=2.3e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1345 $X2=0.1890 $Y2=0.1345
r39 1 25 0.347531 $w=1.965e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1795
+ $Y=0.1345 $X2=0.1785 $Y2=0.1345
r40 9 23 2.44436 $w=1.30368e-07 $l=5e-10 $layer=LIG $thickness=5.22105e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1345
r41 9 25 0.54388 $w=2.16967e-07 $l=1.05119e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1345
r42 9 26 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1345
r43 3 11 1e-05
.ends


*
.SUBCKT AND2x2_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM5@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM5@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND2x2_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1 PM_AND2x2_ASAP7_75t_R%noxref_8
cc_1 N_noxref_8_1 N_MM2_g 0.00242233f
cc_2 N_noxref_8_1 N_NET10_11 0.0371632f
x_PM_AND2x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND2x2_ASAP7_75t_R%noxref_10
cc_3 N_noxref_10_1 N_MM5@2_g 0.00146192f
cc_4 N_noxref_10_1 N_Y_7 0.000839325f
x_PM_AND2x2_ASAP7_75t_R%A VSS A N_MM3_g N_A_1 PM_AND2x2_ASAP7_75t_R%A
cc_5 N_MM3_g N_B_1 0.00148242f
cc_6 N_A N_B_6 0.00192713f
cc_7 N_MM3_g N_MM2_g 0.00784069f
x_PM_AND2x2_ASAP7_75t_R%NET20 VSS N_MM2_s N_MM3_d N_NET20_1
+ PM_AND2x2_ASAP7_75t_R%NET20
cc_8 N_NET20_1 N_MM2_g 0.0173893f
cc_9 N_NET20_1 N_MM3_g 0.0174017f
cc_10 N_NET20_1 N_NET10_11 0.000372959f
x_PM_AND2x2_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_AND2x2_ASAP7_75t_R%noxref_9
cc_11 N_noxref_9_1 N_MM2_g 0.00443199f
cc_12 N_noxref_9_1 N_NET10_12 0.000646344f
cc_13 N_noxref_9_1 N_noxref_8_1 0.00189452f
x_PM_AND2x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND2x2_ASAP7_75t_R%noxref_11
cc_14 N_noxref_11_1 N_MM5@2_g 0.00146434f
cc_15 N_noxref_11_1 N_Y_8 0.000823914f
cc_16 N_noxref_11_1 N_noxref_10_1 0.00178075f
x_PM_AND2x2_ASAP7_75t_R%Y VSS Y N_MM5_d N_MM5@2_d N_MM4_d N_MM4@2_d N_Y_7
+ N_Y_10 N_Y_8 N_Y_15 N_Y_14 N_Y_2 N_Y_1 N_Y_9 PM_AND2x2_ASAP7_75t_R%Y
cc_17 N_Y_7 N_NET10_17 0.000403795f
cc_18 N_Y_7 N_NET10_1 0.00670254f
cc_19 N_Y_10 N_NET10_20 0.000833751f
cc_20 N_Y_8 N_MM5@2_g 0.030884f
cc_21 N_Y_15 N_NET10_21 0.000993501f
cc_22 N_Y_14 N_NET10_19 0.00106582f
cc_23 N_Y_2 N_MM5@2_g 0.00208098f
cc_24 N_Y_1 N_MM5@2_g 0.0021248f
cc_25 N_Y_10 N_NET10_17 0.00304766f
cc_26 N_Y_9 N_NET10_16 0.00318696f
cc_27 N_Y_7 N_MM5_g 0.0370915f
cc_28 N_Y_7 N_MM5@2_g 0.069024f
x_PM_AND2x2_ASAP7_75t_R%B VSS B N_MM2_g N_B_1 N_B_6 N_B_4 N_B_5
+ PM_AND2x2_ASAP7_75t_R%B
x_PM_AND2x2_ASAP7_75t_R%NET10 VSS N_MM5_g N_MM5@2_g N_MM1_d N_MM0_d N_MM2_d
+ N_NET10_18 N_NET10_3 N_NET10_4 N_NET10_13 N_NET10_15 N_NET10_11 N_NET10_12
+ N_NET10_20 N_NET10_14 N_NET10_1 N_NET10_17 N_NET10_16 N_NET10_21 N_NET10_19
+ PM_AND2x2_ASAP7_75t_R%NET10
cc_29 N_NET10_18 N_MM2_g 0.000386915f
cc_30 N_NET10_3 N_B_4 0.000447486f
cc_31 N_NET10_4 N_MM2_g 0.00062799f
cc_32 N_NET10_3 N_B_1 0.000706509f
cc_33 N_NET10_13 N_B_6 0.000809493f
cc_34 N_NET10_15 N_B_5 0.0010232f
cc_35 N_NET10_11 N_B_1 0.00252782f
cc_36 N_NET10_13 N_B_4 0.00365157f
cc_37 N_NET10_12 N_MM2_g 0.0109851f
cc_38 N_NET10_3 N_MM2_g 0.00481441f
cc_39 N_NET10_11 N_MM2_g 0.0507047f
cc_40 N_NET10_13 N_MM3_g 0.000582187f
cc_41 N_NET10_4 N_MM3_g 0.000698578f
cc_42 N_NET10_20 N_A_1 0.000830139f
cc_43 N_NET10_3 N_MM3_g 0.000875883f
cc_44 N_NET10_14 N_A 0.000883808f
cc_45 N_NET10_15 N_A 0.000893673f
cc_46 N_NET10_1 N_A_1 0.00137999f
cc_47 N_NET10_17 N_A 0.00235896f
cc_48 N_NET10_16 N_A 0.00237827f
cc_49 N_NET10_12 N_MM3_g 0.0110241f
cc_50 N_NET10_20 N_A 0.00845511f
cc_51 N_MM5_g N_MM3_g 0.0187013f
*END of AND2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AND2x4_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND2x4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND2x4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND2x4_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0328101f
.ends

.subckt PM_AND2x4_ASAP7_75t_R%NET19 VSS 2 3 1
c1 1 VSS 0.000931474f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AND2x4_ASAP7_75t_R%NET19__2 VSS 2 3 1
c1 1 VSS 0.000911542f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND2x4_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0425255f
.ends

.subckt PM_AND2x4_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0430772f
.ends

.subckt PM_AND2x4_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0430709f
.ends

.subckt PM_AND2x4_ASAP7_75t_R%B VSS 19 3 4 1 5
c1 1 VSS 0.00799663f
c2 3 VSS 0.0361f
c3 4 VSS 0.0360112f
c4 5 VSS 0.00453142f
r1 19 18 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1520 $X2=0.1350 $Y2=0.1477
r2 17 18 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1477
r3 5 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1165 $X2=0.1350 $Y2=0.1350
r4 3 12 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 12 13 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r6 12 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r7 9 13 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r8 8 9 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.1620
+ $Y=0.1350 $X2=0.1475 $Y2=0.1350
r9 7 8 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.1765
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r10 4 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r11 1 7 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r12 1 15 4.63801 $w=1.7681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
r13 4 7 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r14 4 15 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1995 $Y2=0.1350
.ends

.subckt PM_AND2x4_ASAP7_75t_R%A VSS 18 5 6 1 2 7 8 9
c1 1 VSS 0.0041095f
c2 2 VSS 0.00372878f
c3 5 VSS 0.0713176f
c4 6 VSS 0.0820068f
c5 7 VSS 0.0125919f
c6 8 VSS 0.0157395f
c7 9 VSS 0.00566816f
c8 10 VSS 0.00491131f
c9 11 VSS 0.00454475f
r1 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r2 6 2 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1235 $X2=0.2430 $Y2=0.1350
r4 24 25 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0925 $X2=0.2430 $Y2=0.1235
r5 9 23 2.14973 $w=1.32632e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0550 $X2=0.2430 $Y2=0.0455
r6 9 24 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0550 $X2=0.2430 $Y2=0.0925
r7 11 23 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0365 $X2=0.2430 $Y2=0.0455
r8 22 23 4.24844 $w=1.31351e-08 $l=2.83064e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0370 $X2=0.2430 $Y2=0.0455
r9 21 22 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1565
+ $Y=0.0370 $X2=0.2160 $Y2=0.0370
r10 20 21 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1045
+ $Y=0.0370 $X2=0.1565 $Y2=0.0370
r11 8 10 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0920 $Y=0.0370 $X2=0.0810 $Y2=0.0370
r12 8 20 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0920
+ $Y=0.0370 $X2=0.1045 $Y2=0.0370
r13 10 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0370 $X2=0.0810 $Y2=0.0550
r14 18 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1165
r15 15 16 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0730 $X2=0.0810 $Y2=0.0550
r16 7 15 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0945 $X2=0.0810 $Y2=0.0730
r17 7 17 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0945 $X2=0.0810 $Y2=0.1165
r18 5 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r19 18 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AND2x4_ASAP7_75t_R%Y VSS 31 24 25 36 37 44 45 48 49 13 4 18 1 2 16
+ 15 14
c1 1 VSS 0.0102961f
c2 2 VSS 0.0102793f
c3 3 VSS 0.00973187f
c4 4 VSS 0.00974254f
c5 13 VSS 0.00452198f
c6 14 VSS 0.00455497f
c7 15 VSS 0.00443586f
c8 16 VSS 0.00457809f
c9 17 VSS 0.0151256f
c10 18 VSS 0.0137884f
c11 19 VSS 0.00796792f
c12 20 VSS 0.00360644f
c13 21 VSS 0.00355116f
r1 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 4 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r6 2 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r8 44 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r9 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r10 2 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r11 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r12 39 40 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r13 38 39 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r14 18 38 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r15 21 33 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4590 $Y2=0.2125
r16 21 41 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r17 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r18 3 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r19 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r20 36 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r21 32 33 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1740 $X2=0.4590 $Y2=0.2125
r22 31 32 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1740
r23 31 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1340
r24 19 20 9.31081 $w=1.48766e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0830 $X2=0.4590 $Y2=0.0360
r25 19 30 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0830 $X2=0.4590 $Y2=0.1340
r26 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r27 20 29 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r28 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r29 27 28 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r30 26 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r31 17 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r32 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r33 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r34 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r35 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r36 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
.ends

.subckt PM_AND2x4_ASAP7_75t_R%NET9 VSS 12 13 14 15 78 79 82 83 86 87 18 5 4 1
+ 19 3 23 24 26 20 21 17 25 16 28
c1 1 VSS 0.0185201f
c2 3 VSS 0.0108369f
c3 4 VSS 0.00581399f
c4 5 VSS 0.0109141f
c5 12 VSS 0.0814423f
c6 13 VSS 0.081216f
c7 14 VSS 0.0809882f
c8 15 VSS 0.0816609f
c9 16 VSS 0.00569752f
c10 17 VSS 0.00679702f
c11 18 VSS 0.00681187f
c12 19 VSS 0.010186f
c13 20 VSS 0.00163212f
c14 21 VSS 0.00192667f
c15 22 VSS 0.0015419f
c16 23 VSS 0.00381824f
c17 24 VSS 0.0025853f
c18 25 VSS 0.00130469f
c19 26 VSS 0.00129452f
c20 27 VSS 0.00705492f
c21 28 VSS 0.00165958f
r1 87 85 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 3 85 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 17 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 86 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 83 81 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 4 81 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 82 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 79 77 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r10 5 77 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r11 18 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r12 78 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r13 3 75 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1070 $Y2=0.2340
r14 4 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0730
r15 5 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r16 72 73 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1160
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r17 72 75 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1160
+ $Y=0.2340 $X2=0.1070 $Y2=0.2340
r18 71 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r19 70 71 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1615
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r20 19 27 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1795 $Y=0.2340 $X2=0.1890 $Y2=0.2340
r21 19 70 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1795
+ $Y=0.2340 $X2=0.1615 $Y2=0.2340
r22 66 67 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0730 $X2=0.1750 $Y2=0.0730
r23 20 26 0.56619 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1795 $Y=0.0730 $X2=0.1890 $Y2=0.0730
r24 20 67 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1795
+ $Y=0.0730 $X2=0.1750 $Y2=0.0730
r25 62 63 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r26 27 62 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.2025 $Y2=0.2340
r27 26 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0730 $X2=0.1890 $Y2=0.0945
r28 22 25 3.85983 $w=1.51591e-08 $l=2.15058e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2125 $X2=0.1885 $Y2=0.1910
r29 22 27 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2125 $X2=0.1890 $Y2=0.2340
r30 60 61 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1285 $X2=0.1890 $Y2=0.0945
r31 21 25 4.67599 $w=1.48627e-08 $l=2.5005e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1660 $X2=0.1885 $Y2=0.1910
r32 21 60 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1660 $X2=0.1890 $Y2=0.1285
r33 25 59 4.79259 $w=1.48269e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1885 $Y=0.1910 $X2=0.2145 $Y2=0.1910
r34 58 59 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2325
+ $Y=0.1910 $X2=0.2145 $Y2=0.1910
r35 57 58 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1910 $X2=0.2325 $Y2=0.1910
r36 23 28 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1910 $X2=0.2970 $Y2=0.1910
r37 23 57 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1910 $X2=0.2430 $Y2=0.1910
r38 28 53 4.18063 $w=1.6528e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1910 $X2=0.2970 $Y2=0.1660
r39 15 49 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r40 14 43 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r41 13 37 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r42 52 53 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1470 $X2=0.2970 $Y2=0.1660
r43 51 52 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1470
r44 24 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1235 $X2=0.2970 $Y2=0.1350
r45 47 49 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r46 46 47 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r47 44 46 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r48 43 44 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r49 41 43 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r50 40 41 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r51 38 40 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r52 37 38 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r53 35 37 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r54 34 35 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r55 33 34 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r56 31 33 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r57 30 31 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r58 30 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r59 1 30 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r60 1 32 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r61 12 30 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r62 12 32 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r63 12 33 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends


*
.SUBCKT AND2x4_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3@2 N_MM3@2_d N_MM3@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM1@2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@4 N_MM5@4_d N_MM4@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 N_MM5@3_d N_MM4@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@4 N_MM4@4_d N_MM4@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM4@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND2x4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND2x4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND2x4_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND2x4_ASAP7_75t_R%noxref_10
cc_1 N_noxref_10_1 N_MM3@2_g 0.00377658f
cc_2 N_noxref_10_1 N_noxref_9_1 0.00192695f
x_PM_AND2x4_ASAP7_75t_R%NET19 VSS N_MM2_s N_MM3_d N_NET19_1
+ PM_AND2x4_ASAP7_75t_R%NET19
cc_3 N_NET19_1 N_MM0@2_g 0.0174249f
cc_4 N_NET19_1 N_MM1@2_g 0.0174225f
x_PM_AND2x4_ASAP7_75t_R%NET19__2 VSS N_MM3@2_d N_MM2@2_s N_NET19__2_1
+ PM_AND2x4_ASAP7_75t_R%NET19__2
cc_5 N_NET19__2_1 N_MM3@2_g 0.0171391f
cc_6 N_NET19__2_1 N_MM2@2_g 0.0172647f
x_PM_AND2x4_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_AND2x4_ASAP7_75t_R%noxref_9
cc_7 N_noxref_9_1 N_MM3@2_g 0.0018878f
x_PM_AND2x4_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND2x4_ASAP7_75t_R%noxref_11
cc_8 N_noxref_11_1 N_MM4@2_g 0.00148841f
x_PM_AND2x4_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND2x4_ASAP7_75t_R%noxref_12
cc_9 N_noxref_12_1 N_MM4@2_g 0.00148311f
cc_10 N_noxref_12_1 N_noxref_11_1 0.00179123f
x_PM_AND2x4_ASAP7_75t_R%B VSS B N_MM2@2_g N_MM1@2_g N_B_1 N_B_5
+ PM_AND2x4_ASAP7_75t_R%B
cc_11 N_MM2@2_g N_A_1 0.00114338f
cc_12 N_B_1 N_A_2 0.00213481f
cc_13 N_B_5 N_A_7 0.00389092f
cc_14 N_MM1@2_g N_MM0@2_g 0.00717857f
cc_15 N_MM2@2_g N_MM3@2_g 0.00865464f
x_PM_AND2x4_ASAP7_75t_R%A VSS A N_MM3@2_g N_MM0@2_g N_A_1 N_A_2 N_A_7 N_A_8
+ N_A_9 PM_AND2x4_ASAP7_75t_R%A
x_PM_AND2x4_ASAP7_75t_R%Y VSS Y N_MM5_d N_MM5@4_d N_MM5@3_d N_MM5@2_d N_MM4_d
+ N_MM4@4_d N_MM4@3_d N_MM4@2_d N_Y_13 N_Y_4 N_Y_18 N_Y_1 N_Y_2 N_Y_16 N_Y_15
+ N_Y_14 PM_AND2x4_ASAP7_75t_R%Y
cc_16 N_Y_13 N_MM4@3_g 0.000471796f
cc_17 N_Y_13 N_NET9_1 0.00176711f
cc_18 N_Y_13 N_MM4@2_g 0.00349117f
cc_19 N_Y_13 N_NET9_24 0.00108618f
cc_20 N_Y_4 N_MM4@2_g 0.00180894f
cc_21 N_Y_18 N_NET9_28 0.00186061f
cc_22 N_Y_1 N_MM4@4_g 0.00201555f
cc_23 N_Y_2 N_MM4@4_g 0.00226017f
cc_24 N_Y_16 N_NET9_1 0.00973878f
cc_25 N_Y_16 N_MM4@2_g 0.0295521f
cc_26 N_Y_15 N_MM4@4_g 0.0296284f
cc_27 N_Y_14 N_MM4@2_g 0.0659377f
cc_28 N_Y_13 N_MM4_g 0.0364397f
cc_29 N_Y_14 N_MM4@3_g 0.0365158f
cc_30 N_Y_13 N_MM4@4_g 0.0689009f
x_PM_AND2x4_ASAP7_75t_R%NET9 VSS N_MM4_g N_MM4@4_g N_MM4@3_g N_MM4@2_g
+ N_MM1@2_d N_MM0@2_d N_MM2@2_d N_MM2_d N_MM0_d N_MM1_d N_NET9_18 N_NET9_5
+ N_NET9_4 N_NET9_1 N_NET9_19 N_NET9_3 N_NET9_23 N_NET9_24 N_NET9_26 N_NET9_20
+ N_NET9_21 N_NET9_17 N_NET9_25 N_NET9_16 N_NET9_28 PM_AND2x4_ASAP7_75t_R%NET9
cc_31 N_NET9_18 N_MM3@2_g 0.000351058f
cc_32 N_NET9_5 N_MM0@2_g 0.000386029f
cc_33 N_NET9_4 N_A_8 0.00149095f
cc_34 N_NET9_1 N_MM0@2_g 0.000499318f
cc_35 N_NET9_19 N_A_7 0.000612802f
cc_36 N_NET9_3 N_MM3@2_g 0.00072915f
cc_37 N_NET9_1 N_A_2 0.00221358f
cc_38 N_NET9_23 N_A_9 0.00105656f
cc_39 N_NET9_24 N_A_9 0.00106326f
cc_40 N_NET9_26 N_A_8 0.00158403f
cc_41 N_NET9_20 N_A_7 0.002287f
cc_42 N_NET9_18 N_MM0@2_g 0.0109814f
cc_43 N_NET9_21 N_A_9 0.00560086f
cc_44 N_NET9_20 N_A_8 0.00775475f
cc_45 N_MM4_g N_MM0@2_g 0.0172269f
cc_46 N_NET9_17 N_MM3@2_g 0.0267416f
cc_47 N_NET9_17 N_MM1@2_g 0.000358974f
cc_48 N_NET9_5 N_MM1@2_g 0.000395942f
cc_49 N_NET9_25 N_MM1@2_g 0.000439759f
cc_50 N_NET9_4 N_MM1@2_g 0.00307181f
cc_51 N_NET9_3 N_MM2@2_g 0.000724796f
cc_52 N_NET9_20 N_B_5 0.000982047f
cc_53 N_NET9_19 N_B_5 0.00104529f
cc_54 N_NET9_16 N_B_1 0.0036349f
cc_55 N_NET9_18 N_MM1@2_g 0.0109698f
cc_56 N_NET9_17 N_MM2@2_g 0.0110074f
cc_57 N_NET9_21 N_B_5 0.00650067f
cc_58 N_NET9_16 N_MM2@2_g 0.0332658f
cc_59 N_NET9_16 N_MM1@2_g 0.0663395f
*END of AND2x4_ASAP7_75t_R.pxi
.ENDS
** Design:	AND2x6_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND2x6_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND2x6_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND2x6_ASAP7_75t_R%NET19 VSS 2 3 1
c1 1 VSS 0.000931504f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AND2x6_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0425216f
.ends

.subckt PM_AND2x6_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0328146f
.ends

.subckt PM_AND2x6_ASAP7_75t_R%NET19__2 VSS 2 3 1
c1 1 VSS 0.000911348f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND2x6_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0430484f
.ends

.subckt PM_AND2x6_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0430476f
.ends

.subckt PM_AND2x6_ASAP7_75t_R%A VSS 18 5 6 1 2 7 8 9
c1 1 VSS 0.00409969f
c2 2 VSS 0.00365086f
c3 5 VSS 0.0713173f
c4 6 VSS 0.0819871f
c5 7 VSS 0.0124505f
c6 8 VSS 0.0154458f
c7 9 VSS 0.00557908f
c8 10 VSS 0.0048962f
c9 11 VSS 0.00454677f
r1 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r2 6 2 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 25 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1235 $X2=0.2430 $Y2=0.1350
r4 24 25 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0925 $X2=0.2430 $Y2=0.1235
r5 9 23 2.14973 $w=1.32632e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0550 $X2=0.2430 $Y2=0.0455
r6 9 24 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0550 $X2=0.2430 $Y2=0.0925
r7 11 23 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0365 $X2=0.2430 $Y2=0.0455
r8 22 23 4.24844 $w=1.31351e-08 $l=2.83064e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.0370 $X2=0.2430 $Y2=0.0455
r9 21 22 13.8748 $w=1.3e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1565
+ $Y=0.0370 $X2=0.2160 $Y2=0.0370
r10 20 21 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1045
+ $Y=0.0370 $X2=0.1565 $Y2=0.0370
r11 8 10 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0920 $Y=0.0370 $X2=0.0810 $Y2=0.0370
r12 8 20 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0920
+ $Y=0.0370 $X2=0.1045 $Y2=0.0370
r13 10 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0370 $X2=0.0810 $Y2=0.0550
r14 18 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1165
r15 15 16 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0730 $X2=0.0810 $Y2=0.0550
r16 7 15 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0945 $X2=0.0810 $Y2=0.0730
r17 7 17 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0945 $X2=0.0810 $Y2=0.1165
r18 5 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r19 18 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AND2x6_ASAP7_75t_R%B VSS 18 3 4 1 5
c1 1 VSS 0.0081439f
c2 3 VSS 0.0361731f
c3 4 VSS 0.0360924f
c4 5 VSS 0.00469042f
r1 4 14 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 18 17 0.991056 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1520 $X2=0.1350 $Y2=0.1477
r3 16 17 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1477
r4 5 16 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1165 $X2=0.1350 $Y2=0.1350
r5 12 14 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 11 12 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r7 10 11 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r8 8 10 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1475 $Y2=0.1350
r9 7 8 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r10 7 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r11 1 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r12 1 9 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1245 $Y2=0.1350
r13 3 7 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r14 3 9 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1245 $Y2=0.1350
r15 3 10 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
.ends

.subckt PM_AND2x6_ASAP7_75t_R%Y VSS 41 34 35 48 49 58 59 62 63 66 67 70 71 20 2
+ 27 4 5 3 6 26 1 24 23 22 21 19
c1 1 VSS 0.0102319f
c2 2 VSS 0.0101935f
c3 3 VSS 0.00972589f
c4 4 VSS 0.00974227f
c5 5 VSS 0.0107183f
c6 6 VSS 0.0107234f
c7 19 VSS 0.00447365f
c8 20 VSS 0.00435682f
c9 21 VSS 0.00452121f
c10 22 VSS 0.00440531f
c11 23 VSS 0.0043447f
c12 24 VSS 0.00451962f
c13 25 VSS 0.0153355f
c14 26 VSS 0.0136562f
c15 27 VSS 0.00561503f
c16 28 VSS 0.00948619f
c17 29 VSS 0.00966983f
c18 30 VSS 0.00254135f
c19 31 VSS 0.00254135f
r1 71 69 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 6 69 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 24 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 70 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 67 65 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 4 65 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 23 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 66 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r10 2 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r11 22 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r12 62 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r13 6 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r14 4 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r15 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r16 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r17 5 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r18 21 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r19 58 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r20 29 54 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r21 29 31 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4995 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r22 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r23 51 52 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r24 50 51 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r25 26 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r26 5 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r27 31 43 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4590 $Y2=0.2125
r28 31 53 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r29 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r30 3 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r31 20 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r32 48 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r33 28 44 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r34 28 30 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4995 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r35 42 43 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1740 $X2=0.4590 $Y2=0.2125
r36 41 42 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1740
r37 41 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1340
r38 27 30 9.77961 $w=1.39574e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0830 $X2=0.4590 $Y2=0.0360
r39 27 40 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0830 $X2=0.4590 $Y2=0.1340
r40 3 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r41 30 39 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r42 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r43 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r44 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r45 25 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r46 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r47 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r48 1 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r49 19 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r50 34 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
.ends

.subckt PM_AND2x6_ASAP7_75t_R%NET9 VSS 12 13 14 15 16 17 94 95 98 99 102 103 18
+ 20 5 4 1 21 3 25 26 28 22 23 19 27 30
c1 1 VSS 0.0295091f
c2 3 VSS 0.0120611f
c3 4 VSS 0.00703824f
c4 5 VSS 0.0121383f
c5 12 VSS 0.0820544f
c6 13 VSS 0.0818766f
c7 14 VSS 0.0818195f
c8 15 VSS 0.0817733f
c9 16 VSS 0.0816114f
c10 17 VSS 0.0823698f
c11 18 VSS 0.00753415f
c12 19 VSS 0.00863469f
c13 20 VSS 0.00864824f
c14 21 VSS 0.0108007f
c15 22 VSS 0.00224449f
c16 23 VSS 0.00253418f
c17 24 VSS 0.00215482f
c18 25 VSS 0.00442332f
c19 26 VSS 0.0031972f
c20 27 VSS 0.00191681f
c21 28 VSS 0.00190664f
c22 29 VSS 0.00722156f
c23 30 VSS 0.00222908f
r1 103 101 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 3 101 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 19 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 102 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 99 97 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 4 97 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 18 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 98 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 95 93 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r10 5 93 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2160 $X2=0.2305 $Y2=0.2160
r11 20 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2160 $X2=0.2160 $Y2=0.2160
r12 94 20 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2160 $X2=0.2015 $Y2=0.2160
r13 3 91 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1070 $Y2=0.2340
r14 4 82 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0730
r15 5 79 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r16 88 89 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1160
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r17 88 91 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1160
+ $Y=0.2340 $X2=0.1070 $Y2=0.2340
r18 87 89 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r19 86 87 6.17953 $w=1.3e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1615
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r20 21 29 1.03499 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1795 $Y=0.2340 $X2=0.1890 $Y2=0.2340
r21 21 86 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1795
+ $Y=0.2340 $X2=0.1615 $Y2=0.2340
r22 82 83 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0730 $X2=0.1750 $Y2=0.0730
r23 22 28 0.56619 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.1795 $Y=0.0730 $X2=0.1890 $Y2=0.0730
r24 22 83 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1795
+ $Y=0.0730 $X2=0.1750 $Y2=0.0730
r25 78 79 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r26 29 78 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2340 $X2=0.2025 $Y2=0.2340
r27 28 77 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.0730 $X2=0.1890 $Y2=0.0945
r28 24 27 3.85983 $w=1.51591e-08 $l=2.15058e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2125 $X2=0.1885 $Y2=0.1910
r29 24 29 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.2125 $X2=0.1890 $Y2=0.2340
r30 76 77 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1285 $X2=0.1890 $Y2=0.0945
r31 23 27 4.67599 $w=1.48627e-08 $l=2.5005e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1660 $X2=0.1885 $Y2=0.1910
r32 23 76 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1660 $X2=0.1890 $Y2=0.1285
r33 27 75 4.79259 $w=1.48269e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1885 $Y=0.1910 $X2=0.2145 $Y2=0.1910
r34 74 75 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2325
+ $Y=0.1910 $X2=0.2145 $Y2=0.1910
r35 73 74 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1910 $X2=0.2325 $Y2=0.1910
r36 25 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1910 $X2=0.2970 $Y2=0.1910
r37 25 73 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1910 $X2=0.2430 $Y2=0.1910
r38 30 67 4.18063 $w=1.6528e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1910 $X2=0.2970 $Y2=0.1660
r39 17 63 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r40 16 57 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r41 15 51 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r42 14 45 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r43 13 39 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r44 66 67 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1470 $X2=0.2970 $Y2=0.1660
r45 65 66 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1470
r46 26 65 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1235 $X2=0.2970 $Y2=0.1350
r47 61 63 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r48 60 61 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r49 58 60 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r50 57 58 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r51 55 57 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r52 54 55 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r53 52 54 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r54 51 52 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r55 49 51 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r56 48 49 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r57 46 48 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r58 45 46 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r59 43 45 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r60 42 43 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r61 40 42 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r62 39 40 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r63 37 39 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r64 36 37 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r65 35 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r66 33 35 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r67 32 33 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r68 32 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r69 1 32 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r70 1 34 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r71 12 32 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r72 12 34 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r73 12 35 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends


*
.SUBCKT AND2x6_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3@2 N_MM3@2_d N_MM3@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM1_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM1@2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@6 N_MM5@6_d N_MM4@6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@5 N_MM5@5_d N_MM4@5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@4 N_MM5@4_d N_MM4@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 N_MM5@3_d N_MM4@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM4@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 N_MM1@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@6 N_MM4@6_d N_MM4@6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@5 N_MM4@5_d N_MM4@5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@4 N_MM4@4_d N_MM4@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@3 N_MM4@3_d N_MM4@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND2x6_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND2x6_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND2x6_ASAP7_75t_R%NET19 VSS N_MM2_s N_MM3_d N_NET19_1
+ PM_AND2x6_ASAP7_75t_R%NET19
cc_1 N_NET19_1 N_MM0@2_g 0.0174243f
cc_2 N_NET19_1 N_MM1@2_g 0.0174231f
x_PM_AND2x6_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_AND2x6_ASAP7_75t_R%noxref_9
cc_3 N_noxref_9_1 N_MM3@2_g 0.0018875f
x_PM_AND2x6_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND2x6_ASAP7_75t_R%noxref_10
cc_4 N_noxref_10_1 N_MM3@2_g 0.00377863f
cc_5 N_noxref_10_1 N_noxref_9_1 0.00192606f
x_PM_AND2x6_ASAP7_75t_R%NET19__2 VSS N_MM3@2_d N_MM2@2_s N_NET19__2_1
+ PM_AND2x6_ASAP7_75t_R%NET19__2
cc_6 N_NET19__2_1 N_MM3@2_g 0.0171375f
cc_7 N_NET19__2_1 N_MM1_g 0.0172664f
x_PM_AND2x6_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND2x6_ASAP7_75t_R%noxref_11
cc_8 N_noxref_11_1 N_MM4@2_g 0.00150354f
x_PM_AND2x6_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND2x6_ASAP7_75t_R%noxref_12
cc_9 N_noxref_12_1 N_MM4@2_g 0.0014998f
cc_10 N_noxref_12_1 N_noxref_11_1 0.00179873f
x_PM_AND2x6_ASAP7_75t_R%A VSS A N_MM3@2_g N_MM0@2_g N_A_1 N_A_2 N_A_7 N_A_8
+ N_A_9 PM_AND2x6_ASAP7_75t_R%A
x_PM_AND2x6_ASAP7_75t_R%B VSS B N_MM1_g N_MM1@2_g N_B_1 N_B_5
+ PM_AND2x6_ASAP7_75t_R%B
cc_11 N_MM1_g N_A_1 0.00114338f
cc_12 N_B_1 N_A_2 0.0021047f
cc_13 N_B_5 N_A_7 0.00409874f
cc_14 N_MM1@2_g N_MM0@2_g 0.00717857f
cc_15 N_MM1_g N_MM3@2_g 0.00865846f
x_PM_AND2x6_ASAP7_75t_R%Y VSS Y N_MM5_d N_MM5@6_d N_MM5@5_d N_MM5@4_d N_MM5@3_d
+ N_MM5@2_d N_MM4_d N_MM4@6_d N_MM4@5_d N_MM4@4_d N_MM4@3_d N_MM4@2_d N_Y_20
+ N_Y_2 N_Y_27 N_Y_4 N_Y_5 N_Y_3 N_Y_6 N_Y_26 N_Y_1 N_Y_24 N_Y_23 N_Y_22 N_Y_21
+ N_Y_19 PM_AND2x6_ASAP7_75t_R%Y
cc_16 N_Y_20 N_NET9_25 0.000430233f
cc_17 N_Y_20 N_MM4@5_g 0.0368092f
cc_18 N_Y_20 N_NET9_1 0.000509989f
cc_19 N_Y_20 N_MM4@2_g 0.00172235f
cc_20 N_Y_20 N_MM4@6_g 0.00172386f
cc_21 N_Y_2 N_NET9_26 0.00109265f
cc_22 N_Y_27 N_NET9_1 0.00164462f
cc_23 N_Y_4 N_MM4@4_g 0.00171563f
cc_24 N_Y_5 N_MM4@2_g 0.00175132f
cc_25 N_Y_3 N_MM4@4_g 0.00177046f
cc_26 N_Y_6 N_MM4@2_g 0.00178578f
cc_27 N_Y_26 N_NET9_30 0.00187952f
cc_28 N_Y_1 N_MM4@6_g 0.00199191f
cc_29 N_Y_2 N_MM4@6_g 0.00238411f
cc_30 N_Y_24 N_MM4@2_g 0.0293154f
cc_31 N_Y_23 N_MM4@4_g 0.0293657f
cc_32 N_Y_22 N_MM4@6_g 0.0295237f
cc_33 N_Y_23 N_NET9_1 0.0148994f
cc_34 N_Y_21 N_MM4@2_g 0.0655025f
cc_35 N_Y_19 N_MM4@6_g 0.0657214f
cc_36 N_Y_19 N_MM4_g 0.0362284f
cc_37 N_Y_21 N_MM4@3_g 0.0363028f
cc_38 N_Y_20 N_MM4@4_g 0.068571f
x_PM_AND2x6_ASAP7_75t_R%NET9 VSS N_MM4_g N_MM4@6_g N_MM4@5_g N_MM4@4_g
+ N_MM4@3_g N_MM4@2_g N_MM1@2_d N_MM0@2_d N_MM2@2_d N_MM2_d N_MM0_d N_MM1_d
+ N_NET9_18 N_NET9_20 N_NET9_5 N_NET9_4 N_NET9_1 N_NET9_21 N_NET9_3 N_NET9_25
+ N_NET9_26 N_NET9_28 N_NET9_22 N_NET9_23 N_NET9_19 N_NET9_27 N_NET9_30
+ PM_AND2x6_ASAP7_75t_R%NET9
cc_39 N_NET9_18 N_MM3@2_g 0.000248936f
cc_40 N_NET9_20 N_MM3@2_g 0.000351058f
cc_41 N_NET9_5 N_MM0@2_g 0.000386029f
cc_42 N_NET9_4 N_A_8 0.00149095f
cc_43 N_NET9_1 N_MM0@2_g 0.000457863f
cc_44 N_NET9_21 N_A_7 0.000612742f
cc_45 N_NET9_3 N_MM3@2_g 0.00072915f
cc_46 N_NET9_1 N_A_2 0.00213997f
cc_47 N_NET9_25 N_A_9 0.00102348f
cc_48 N_NET9_26 N_A_9 0.00106321f
cc_49 N_NET9_28 N_A_8 0.00158403f
cc_50 N_NET9_22 N_A_7 0.00228385f
cc_51 N_NET9_20 N_MM0@2_g 0.0109814f
cc_52 N_NET9_23 N_A_9 0.00569321f
cc_53 N_NET9_22 N_A_8 0.00751753f
cc_54 N_MM4_g N_MM0@2_g 0.0172269f
cc_55 N_NET9_19 N_MM3@2_g 0.0264852f
cc_56 N_NET9_20 N_MM1@2_g 0.0113276f
cc_57 N_NET9_19 N_MM1@2_g 0.000358974f
cc_58 N_NET9_5 N_MM1@2_g 0.000395942f
cc_59 N_NET9_27 N_MM1@2_g 0.000439759f
cc_60 N_NET9_4 N_MM1@2_g 0.00307181f
cc_61 N_NET9_3 N_MM1_g 0.000724796f
cc_62 N_NET9_22 N_B_5 0.000982027f
cc_63 N_NET9_21 N_B_5 0.00104526f
cc_64 N_NET9_18 N_B_1 0.0036349f
cc_65 N_NET9_19 N_MM1_g 0.0110074f
cc_66 N_NET9_23 N_B_5 0.00661767f
cc_67 N_NET9_18 N_MM1_g 0.0332658f
cc_68 N_NET9_18 N_MM1@2_g 0.0659993f
*END of AND2x6_ASAP7_75t_R.pxi
.ENDS
** Design:	AND3x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND3x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND3x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND3x1_ASAP7_75t_R%NET72 VSS 2 3 1
c1 1 VSS 0.000987086f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND3x1_ASAP7_75t_R%NET71 VSS 2 3 1
c1 1 VSS 0.000946636f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AND3x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00475895f
.ends

.subckt PM_AND3x1_ASAP7_75t_R%C VSS 4 3 1
c1 1 VSS 0.00609658f
c2 3 VSS 0.0832568f
c3 4 VSS 0.0044226f
r1 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AND3x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00502011f
.ends

.subckt PM_AND3x1_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00295585f
c2 3 VSS 0.0430375f
c3 4 VSS 0.0123056f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AND3x1_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.0055202f
c2 3 VSS 0.0460541f
c3 4 VSS 0.00419919f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AND3x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00478072f
.ends

.subckt PM_AND3x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00485512f
.ends

.subckt PM_AND3x1_ASAP7_75t_R%Y VSS 23 15 30 7 12 2 9 1 8 11 10
c1 1 VSS 0.00726004f
c2 2 VSS 0.0069828f
c3 7 VSS 0.00362691f
c4 8 VSS 0.00357137f
c5 9 VSS 0.00265558f
c6 10 VSS 0.00124923f
c7 11 VSS 0.00158019f
c8 12 VSS 0.00280561f
c9 13 VSS 0.000875084f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2150
r4 26 27 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2035 $X2=0.2700 $Y2=0.2150
r5 12 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1920 $X2=0.2835 $Y2=0.1920
r6 12 26 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1920 $X2=0.2700 $Y2=0.2035
r7 13 24 4.99922 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1920 $X2=0.2970 $Y2=0.1655
r8 13 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1920 $X2=0.2835 $Y2=0.1920
r9 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1655
r10 23 22 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1455
r11 21 22 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1455
r12 10 20 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1100 $X2=0.2970 $Y2=0.0850
r13 10 21 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1100 $X2=0.2970 $Y2=0.1350
r14 19 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0850 $X2=0.2970 $Y2=0.0850
r15 18 19 1.86571 $w=1.62e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2710 $Y=0.0850 $X2=0.2835 $Y2=0.0850
r16 11 17 2.31735 $w=1.34762e-08 $l=2.01556e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2620 $Y=0.0850 $X2=0.2700 $Y2=0.0665
r17 11 18 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2620
+ $Y=0.0850 $X2=0.2710 $Y2=0.0850
r18 16 17 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0480 $X2=0.2700 $Y2=0.0665
r19 9 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0365 $X2=0.2700 $Y2=0.0480
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0480
r21 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r22 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_AND3x1_ASAP7_75t_R%NET61 VSS 12 57 60 61 63 4 17 16 14 3 13 5 15 21
+ 19 18 20 22 1
c1 1 VSS 0.00355272f
c2 3 VSS 0.00633995f
c3 4 VSS 0.00848461f
c4 5 VSS 0.00984761f
c5 12 VSS 0.0805186f
c6 13 VSS 0.00297077f
c7 14 VSS 0.00390004f
c8 15 VSS 0.0049272f
c9 16 VSS 0.01774f
c10 17 VSS 0.0168878f
c11 18 VSS 0.00216304f
c12 19 VSS 0.00215265f
c13 20 VSS 0.00313816f
c14 21 VSS 0.000410321f
c15 22 VSS 0.00249594f
r1 63 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 14 62 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 5 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 15 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 60 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 57 56 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r8 13 56 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r9 4 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r10 5 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r11 3 44 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r12 54 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 52 55 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 51 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r17 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 47 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r19 46 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r20 17 22 2.60893 $w=1.47857e-08 $l=1.84391e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2070 $Y=0.2340 $X2=0.2250 $Y2=0.2300
r21 17 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r22 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r23 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r24 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r25 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r26 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r27 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r28 16 20 2.65995 $w=1.48966e-08 $l=1.83371e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2070 $Y=0.0360 $X2=0.2250 $Y2=0.0395
r29 16 38 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 22 35 3.42509 $w=1.44286e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.2300 $X2=0.2250 $Y2=0.2125
r31 20 33 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0395 $X2=0.2250 $Y2=0.0575
r32 34 35 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1915 $X2=0.2250 $Y2=0.2125
r33 19 21 5.4656 $w=1.45789e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1635 $X2=0.2250 $Y2=0.1350
r34 19 34 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1635 $X2=0.2250 $Y2=0.1915
r35 32 33 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0730 $X2=0.2250 $Y2=0.0575
r36 31 32 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0850 $X2=0.2250 $Y2=0.0730
r37 18 21 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1100 $X2=0.2250 $Y2=0.1350
r38 18 31 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1100 $X2=0.2250 $Y2=0.0850
r39 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2365
+ $Y=0.1350 $X2=0.2480 $Y2=0.1350
r40 21 27 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1350 $X2=0.2365 $Y2=0.1350
r41 12 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r42 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2480 $Y2=0.1350
r43 4 14 1e-05
r44 3 13 1e-05
.ends


*
.SUBCKT AND3x1_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND3x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND3x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND3x1_ASAP7_75t_R%NET72 VSS N_MM0_s N_MM1_d N_NET72_1
+ PM_AND3x1_ASAP7_75t_R%NET72
cc_1 N_NET72_1 N_MM0_g 0.0173834f
cc_2 N_NET72_1 N_MM1_g 0.0173268f
x_PM_AND3x1_ASAP7_75t_R%NET71 VSS N_MM1_s N_MM2_d N_NET71_1
+ PM_AND3x1_ASAP7_75t_R%NET71
cc_3 N_NET71_1 N_MM1_g 0.0173618f
cc_4 N_NET71_1 N_MM2_g 0.0172341f
x_PM_AND3x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND3x1_ASAP7_75t_R%noxref_11
cc_5 N_noxref_11_1 N_MM0_g 0.00163416f
cc_6 N_noxref_11_1 N_NET61_14 0.0381679f
cc_7 N_noxref_11_1 N_noxref_10_1 0.00179524f
x_PM_AND3x1_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 PM_AND3x1_ASAP7_75t_R%C
cc_8 N_MM2_g N_B_1 0.00111472f
cc_9 N_C N_B_4 0.00487848f
cc_10 N_MM2_g N_MM1_g 0.00620376f
x_PM_AND3x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND3x1_ASAP7_75t_R%noxref_10
cc_11 N_noxref_10_1 N_MM0_g 0.00163963f
cc_12 N_noxref_10_1 N_NET61_13 0.0379029f
x_PM_AND3x1_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_AND3x1_ASAP7_75t_R%A
x_PM_AND3x1_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4 PM_AND3x1_ASAP7_75t_R%B
cc_13 N_B_1 N_A_1 0.00124528f
cc_14 N_B_4 N_A_4 0.00470481f
cc_15 N_MM1_g N_MM0_g 0.00631197f
x_PM_AND3x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AND3x1_ASAP7_75t_R%noxref_13
cc_16 N_noxref_13_1 N_MM7_g 0.0015058f
cc_17 N_noxref_13_1 N_Y_8 0.0383802f
cc_18 N_noxref_13_1 N_noxref_12_1 0.00177124f
x_PM_AND3x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND3x1_ASAP7_75t_R%noxref_12
cc_19 N_noxref_12_1 N_MM7_g 0.00150004f
cc_20 N_noxref_12_1 N_Y_7 0.0383247f
x_PM_AND3x1_ASAP7_75t_R%Y VSS Y N_MM7_d N_MM6_d N_Y_7 N_Y_12 N_Y_2 N_Y_9 N_Y_1
+ N_Y_8 N_Y_11 N_Y_10 PM_AND3x1_ASAP7_75t_R%Y
cc_21 N_Y_7 N_NET61_19 0.000364824f
cc_22 N_Y_7 N_NET61_21 0.000366047f
cc_23 N_Y_7 N_NET61_20 0.000487927f
cc_24 N_Y_12 N_NET61_22 0.000526774f
cc_25 N_Y_2 N_NET61_1 0.000932265f
cc_26 N_Y_9 N_NET61_18 0.00107273f
cc_27 N_Y_1 N_MM7_g 0.00143217f
cc_28 N_Y_2 N_MM7_g 0.00146079f
cc_29 N_Y_8 N_NET61_1 0.00253602f
cc_30 N_Y_11 N_NET61_18 0.00277735f
cc_31 N_Y_10 N_NET61_21 0.00305927f
cc_32 N_Y_12 N_NET61_19 0.00366719f
cc_33 N_Y_8 N_MM7_g 0.015204f
cc_34 N_Y_7 N_MM7_g 0.0549648f
x_PM_AND3x1_ASAP7_75t_R%NET61 VSS N_MM7_g N_MM0_d N_MM4_d N_MM5_d N_MM3_d
+ N_NET61_4 N_NET61_17 N_NET61_16 N_NET61_14 N_NET61_3 N_NET61_13 N_NET61_5
+ N_NET61_15 N_NET61_21 N_NET61_19 N_NET61_18 N_NET61_20 N_NET61_22 N_NET61_1
+ PM_AND3x1_ASAP7_75t_R%NET61
cc_35 N_NET61_4 N_A_1 0.000806868f
cc_36 N_NET61_17 N_A_4 0.00127592f
cc_37 N_NET61_16 N_A_4 0.00139765f
cc_38 N_NET61_4 N_MM0_g 0.00149842f
cc_39 N_NET61_14 N_A_1 0.00171038f
cc_40 N_NET61_3 N_MM0_g 0.00185225f
cc_41 N_NET61_4 N_A_4 0.00423857f
cc_42 N_NET61_14 N_MM0_g 0.0154757f
cc_43 N_NET61_13 N_MM0_g 0.055319f
cc_44 N_NET61_5 N_MM1_g 0.00156774f
cc_45 N_NET61_15 N_B_1 0.000695851f
cc_46 N_NET61_17 N_B_4 0.00116703f
cc_47 N_NET61_16 N_B_4 0.00144788f
cc_48 N_NET61_5 N_B_4 0.0033365f
cc_49 N_NET61_15 N_MM1_g 0.0360616f
cc_50 N_NET61_21 N_MM2_g 0.00084602f
cc_51 N_NET61_17 N_MM2_g 0.000886464f
cc_52 N_NET61_15 N_C_1 0.000932477f
cc_53 N_NET61_16 N_C 0.0010537f
cc_54 N_NET61_5 N_MM2_g 0.00118598f
cc_55 N_MM7_g N_MM2_g 0.00164643f
cc_56 N_NET61_19 N_C 0.00234074f
cc_57 N_NET61_18 N_C 0.00236963f
cc_58 N_NET61_21 N_C 0.00862319f
cc_59 N_NET61_15 N_MM2_g 0.0372324f
*END of AND3x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AND3x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND3x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND3x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND3x2_ASAP7_75t_R%NET72 VSS 2 3 1
c1 1 VSS 0.0009878f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND3x2_ASAP7_75t_R%NET71 VSS 2 3 1
c1 1 VSS 0.00096146f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AND3x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00491954f
.ends

.subckt PM_AND3x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0423674f
.ends

.subckt PM_AND3x2_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00514754f
c2 3 VSS 0.0459051f
c3 4 VSS 0.00388592f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AND3x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0423639f
.ends

.subckt PM_AND3x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00481838f
.ends

.subckt PM_AND3x2_ASAP7_75t_R%C VSS 8 3 4 1
c1 1 VSS 0.00628382f
c2 3 VSS 0.0831145f
c3 4 VSS 0.00421277f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AND3x2_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00295877f
c2 3 VSS 0.0430144f
c3 4 VSS 0.0123358f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AND3x2_ASAP7_75t_R%Y VSS 28 20 21 36 37 7 2 15 13 14 10 1 9 8
c1 1 VSS 0.00849243f
c2 2 VSS 0.0084707f
c3 7 VSS 0.00460385f
c4 8 VSS 0.00453308f
c5 9 VSS 0.000968163f
c6 10 VSS 0.00122802f
c7 11 VSS 0.00670742f
c8 12 VSS 0.0066262f
c9 13 VSS 0.00726087f
c10 14 VSS 0.00251346f
c11 15 VSS 0.00310057f
c12 16 VSS 0.00348648f
c13 17 VSS 0.00348648f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 36 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r6 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2700 $Y2=0.2160
r7 10 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1865 $X2=0.2700 $Y2=0.1980
r8 15 31 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2815 $Y2=0.2340
r9 15 33 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2700 $Y2=0.2160
r10 12 17 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3130 $Y=0.2340 $X2=0.3510 $Y2=0.2340
r11 12 31 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.2340 $X2=0.2815 $Y2=0.2340
r12 17 30 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.2045
r13 29 30 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1660 $X2=0.3510 $Y2=0.2045
r14 28 29 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1475 $X2=0.3510 $Y2=0.1660
r15 28 27 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1475 $X2=0.3510 $Y2=0.1455
r16 26 27 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1455
r17 25 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1060 $X2=0.3510 $Y2=0.1350
r18 13 16 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0655 $X2=0.3510 $Y2=0.0360
r19 13 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0655 $X2=0.3510 $Y2=0.1060
r20 16 24 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0360 $X2=0.3130 $Y2=0.0360
r21 11 14 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2815 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r22 11 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2815
+ $Y=0.0360 $X2=0.3130 $Y2=0.0360
r23 9 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0720
r24 9 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0360
r25 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0720
r26 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r27 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r28 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r29 20 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_AND3x2_ASAP7_75t_R%NET61 VSS 12 13 59 62 63 65 15 4 18 17 14 3 5 16
+ 1 23 20 19 24 21 22
c1 1 VSS 0.00680619f
c2 3 VSS 0.00714173f
c3 4 VSS 0.0093199f
c4 5 VSS 0.009929f
c5 12 VSS 0.0807439f
c6 13 VSS 0.0808977f
c7 14 VSS 0.00487218f
c8 15 VSS 0.00582581f
c9 16 VSS 0.00662903f
c10 17 VSS 0.0192795f
c11 18 VSS 0.0189775f
c12 19 VSS 0.00260024f
c13 20 VSS 0.00254365f
c14 21 VSS 0.00114514f
c15 22 VSS 0.00286631f
c16 23 VSS 0.000171908f
c17 24 VSS 0.00294571f
r1 65 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 15 64 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r4 5 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r5 16 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r6 62 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r7 59 58 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r8 14 58 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r9 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r10 5 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r11 3 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r12 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 54 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r17 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 49 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r19 48 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r20 18 24 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.2340 $X2=0.2250 $Y2=0.2340
r21 18 48 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r22 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r23 44 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r24 43 44 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r25 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r26 41 42 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r27 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r28 17 22 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.0360 $X2=0.2250 $Y2=0.0360
r29 17 40 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 24 39 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.2340 $X2=0.2250 $Y2=0.2125
r31 22 37 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0360 $X2=0.2250 $Y2=0.0575
r32 38 39 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1920 $X2=0.2250 $Y2=0.2125
r33 20 23 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1640 $X2=0.2250 $Y2=0.1350
r34 20 38 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1640 $X2=0.2250 $Y2=0.1920
r35 36 37 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0780 $X2=0.2250 $Y2=0.0575
r36 19 23 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1060 $X2=0.2250 $Y2=0.1350
r37 19 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1060 $X2=0.2250 $Y2=0.0780
r38 23 33 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1350 $X2=0.2475 $Y2=0.1350
r39 13 31 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r40 21 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2700 $Y=0.1350
+ $X2=0.2700 $Y2=0.1350
r41 21 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2475 $Y2=0.1350
r42 29 31 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r43 28 29 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r44 27 28 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r45 12 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r46 1 26 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r47 1 27 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r48 12 26 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r49 12 27 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r50 4 15 1e-05
r51 3 14 1e-05
.ends


*
.SUBCKT AND3x2_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM7@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM7@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND3x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND3x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND3x2_ASAP7_75t_R%NET72 VSS N_MM0_s N_MM1_d N_NET72_1
+ PM_AND3x2_ASAP7_75t_R%NET72
cc_1 N_NET72_1 N_MM0_g 0.0172784f
cc_2 N_NET72_1 N_MM1_g 0.0174316f
x_PM_AND3x2_ASAP7_75t_R%NET71 VSS N_MM1_s N_MM2_d N_NET71_1
+ PM_AND3x2_ASAP7_75t_R%NET71
cc_3 N_NET71_1 N_MM1_g 0.0173366f
cc_4 N_NET71_1 N_MM2_g 0.017371f
x_PM_AND3x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND3x2_ASAP7_75t_R%noxref_10
cc_5 N_noxref_10_1 N_MM0_g 0.00164127f
cc_6 N_noxref_10_1 N_NET61_3 0.000544435f
cc_7 N_noxref_10_1 N_NET61_14 0.037465f
x_PM_AND3x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND3x2_ASAP7_75t_R%noxref_12
cc_8 N_noxref_12_1 N_MM7@2_g 0.00148611f
cc_9 N_noxref_12_1 N_Y_7 0.000838993f
x_PM_AND3x2_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4 PM_AND3x2_ASAP7_75t_R%B
cc_10 N_B_1 N_A_1 0.00119868f
cc_11 N_B_4 N_A_4 0.00482971f
cc_12 N_MM1_g N_MM0_g 0.00632357f
x_PM_AND3x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AND3x2_ASAP7_75t_R%noxref_13
cc_13 N_noxref_13_1 N_MM7@2_g 0.00148173f
cc_14 N_noxref_13_1 N_Y_8 0.000837332f
cc_15 N_noxref_13_1 N_noxref_12_1 0.00178044f
x_PM_AND3x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND3x2_ASAP7_75t_R%noxref_11
cc_16 N_noxref_11_1 N_MM0_g 0.00163109f
cc_17 N_noxref_11_1 N_NET61_4 0.000542785f
cc_18 N_noxref_11_1 N_NET61_15 0.0375734f
cc_19 N_noxref_11_1 N_noxref_10_1 0.00179327f
x_PM_AND3x2_ASAP7_75t_R%C VSS C N_MM2_g N_C_4 N_C_1 PM_AND3x2_ASAP7_75t_R%C
cc_20 N_MM2_g N_B_1 0.00111958f
cc_21 N_C_4 N_B_4 0.00471089f
cc_22 N_MM2_g N_MM1_g 0.00621528f
x_PM_AND3x2_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_AND3x2_ASAP7_75t_R%A
x_PM_AND3x2_ASAP7_75t_R%Y VSS Y N_MM7_d N_MM7@2_d N_MM6_d N_MM6@2_d N_Y_7 N_Y_2
+ N_Y_15 N_Y_13 N_Y_14 N_Y_10 N_Y_1 N_Y_9 N_Y_8 PM_AND3x2_ASAP7_75t_R%Y
cc_23 N_Y_7 N_NET61_19 0.00042797f
cc_24 N_Y_7 N_NET61_20 0.000434958f
cc_25 N_Y_2 N_NET61_1 0.000934643f
cc_26 N_Y_15 N_NET61_24 0.00108555f
cc_27 N_Y_13 N_NET61_21 0.00108569f
cc_28 N_Y_14 N_NET61_22 0.0011045f
cc_29 N_Y_10 N_NET61_21 0.00162287f
cc_30 N_Y_1 N_MM7@2_g 0.00201685f
cc_31 N_Y_2 N_MM7@2_g 0.00213926f
cc_32 N_Y_10 N_NET61_20 0.00310566f
cc_33 N_Y_9 N_NET61_19 0.0031837f
cc_34 N_Y_8 N_NET61_1 0.00430298f
cc_35 N_Y_8 N_MM7@2_g 0.0299229f
cc_36 N_Y_7 N_MM7_g 0.0372873f
cc_37 N_Y_7 N_MM7@2_g 0.0696394f
x_PM_AND3x2_ASAP7_75t_R%NET61 VSS N_MM7_g N_MM7@2_g N_MM0_d N_MM4_d N_MM5_d
+ N_MM3_d N_NET61_15 N_NET61_4 N_NET61_18 N_NET61_17 N_NET61_14 N_NET61_3
+ N_NET61_5 N_NET61_16 N_NET61_1 N_NET61_23 N_NET61_20 N_NET61_19 N_NET61_24
+ N_NET61_21 N_NET61_22 PM_AND3x2_ASAP7_75t_R%NET61
cc_38 N_NET61_15 N_MM0_g 0.0158982f
cc_39 N_NET61_4 N_A_1 0.000796061f
cc_40 N_NET61_18 N_A_4 0.00125745f
cc_41 N_NET61_17 N_A_4 0.00139159f
cc_42 N_NET61_4 N_MM0_g 0.00150047f
cc_43 N_NET61_14 N_A_1 0.00176798f
cc_44 N_NET61_3 N_MM0_g 0.00186169f
cc_45 N_NET61_4 N_A_4 0.00410008f
cc_46 N_NET61_14 N_MM0_g 0.0550147f
cc_47 N_NET61_3 N_MM1_g 0.000290107f
cc_48 N_NET61_5 N_MM1_g 0.00155097f
cc_49 N_NET61_16 N_B_1 0.000671689f
cc_50 N_NET61_18 N_B_4 0.0011541f
cc_51 N_NET61_17 N_B_4 0.00145187f
cc_52 N_NET61_5 N_B_4 0.00319745f
cc_53 N_NET61_16 N_MM1_g 0.035786f
cc_54 N_NET61_1 N_MM2_g 0.000502485f
cc_55 N_NET61_23 N_MM2_g 0.000745876f
cc_56 N_NET61_18 N_C_4 0.000860466f
cc_57 N_NET61_16 N_C_1 0.000978972f
cc_58 N_NET61_17 N_C_4 0.00104319f
cc_59 N_NET61_5 N_MM2_g 0.00117549f
cc_60 N_MM7_g N_MM2_g 0.0016304f
cc_61 N_NET61_20 N_C_4 0.00230531f
cc_62 N_NET61_19 N_C_4 0.00235793f
cc_63 N_NET61_23 N_C_4 0.00768959f
cc_64 N_NET61_16 N_MM2_g 0.0368961f
*END of AND3x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AND3x4_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND3x4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND3x4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND3x4_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0421167f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00654073f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.04232f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0422729f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%NET90 VSS 11 14 23 26 9 7 1 2 8
c1 1 VSS 0.00994822f
c2 2 VSS 0.00478523f
c3 7 VSS 0.00457148f
c4 8 VSS 0.00225287f
c5 9 VSS 0.0233045f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r2 24 25 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5500 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r3 2 24 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5380 $Y=0.0675 $X2=0.5500 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5380 $Y2=0.0675
r5 23 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r6 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r7 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5015
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r8 18 19 19.9377 $w=1.3e-08 $l=8.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.0360 $X2=0.5015 $Y2=0.0360
r9 17 18 15.1573 $w=1.3e-08 $l=6.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.4160 $Y2=0.0360
r10 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r11 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r12 9 15 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r13 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r14 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r15 12 13 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r16 1 12 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0675 $X2=0.3340 $Y2=0.0675
r17 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r18 11 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00575838f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%B VSS 18 3 4 5 1 7 6
c1 1 VSS 0.0124845f
c2 3 VSS 0.0460733f
c3 4 VSS 0.0474859f
c4 5 VSS 0.00501515f
c5 6 VSS 0.00398287f
c6 7 VSS 0.00497751f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1980 $X2=0.5130 $Y2=0.1665
r2 4 16 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 18 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1665
r4 18 5 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1215
r5 5 6 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1215 $X2=0.5130 $Y2=0.1080
r6 14 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r7 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r8 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r9 10 12 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.5225 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r10 9 10 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5225 $Y2=0.1350
r11 18 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r12 1 9 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r13 1 11 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.5035
+ $Y=0.1350 $X2=0.5025 $Y2=0.1350
r14 3 9 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r15 3 11 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5025 $Y2=0.1350
r16 3 12 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00485514f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.041883f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00620128f
.ends

.subckt PM_AND3x4_ASAP7_75t_R%C VSS 19 3 4 5 1
c1 1 VSS 0.0118327f
c2 3 VSS 0.0839083f
c3 4 VSS 0.0475066f
c4 5 VSS 0.00695663f
r1 19 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1215
r2 5 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1080 $X2=0.3510 $Y2=0.1215
r3 4 13 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r4 19 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r5 12 13 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 10 12 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3415 $Y2=0.1350
r7 9 10 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.3240
+ $Y=0.1350 $X2=0.3385 $Y2=0.1350
r8 8 9 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.3095
+ $Y=0.1350 $X2=0.3240 $Y2=0.1350
r9 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r10 1 7 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r11 1 8 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r12 3 7 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r13 3 8 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends

.subckt PM_AND3x4_ASAP7_75t_R%A VSS 18 3 4 5 1 7 6
c1 1 VSS 0.00867277f
c2 3 VSS 0.00894989f
c3 4 VSS 0.0457788f
c4 5 VSS 0.00417405f
c5 6 VSS 0.00368975f
c6 7 VSS 0.00405322f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1980 $X2=0.6210 $Y2=0.1665
r2 18 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1665
r3 18 5 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1215
r4 5 6 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1215 $X2=0.6210 $Y2=0.1080
r5 3 14 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r6 14 15 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6305 $Y2=0.1350
r7 18 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
r8 11 15 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6305 $Y2=0.1350
r9 10 11 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6335 $Y2=0.1350
r10 9 10 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r11 4 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r12 1 9 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r13 1 17 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6855 $Y2=0.1350
r14 4 9 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r15 4 17 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.6750 $Y=0.1350 $X2=0.6855 $Y2=0.1350
.ends

.subckt PM_AND3x4_ASAP7_75t_R%Y VSS 33 24 25 37 38 46 47 50 51 13 4 15 16 14 19
+ 18 2 1 3
c1 1 VSS 0.00991592f
c2 2 VSS 0.0100045f
c3 3 VSS 0.0102305f
c4 4 VSS 0.010175f
c5 13 VSS 0.0043894f
c6 14 VSS 0.00453751f
c7 15 VSS 0.00441579f
c8 16 VSS 0.0045108f
c9 17 VSS 0.00740825f
c10 18 VSS 0.0199078f
c11 19 VSS 0.0190772f
c12 20 VSS 0.00328496f
c13 21 VSS 0.00335265f
r1 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 4 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 50 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 47 45 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r6 2 45 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r7 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r8 46 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r9 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2125 $Y2=0.2340
r10 2 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r11 40 41 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.2125 $Y2=0.2340
r12 39 40 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r13 19 39 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r14 19 21 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r15 21 34 9.544 $w=1.48375e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.1860
r16 38 36 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r17 3 36 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r18 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r19 37 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r20 33 34 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1465 $X2=0.0270 $Y2=0.1860
r21 33 32 0.349785 $w=1.3e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1465 $X2=0.0270 $Y2=0.1450
r22 31 32 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1450
r23 17 20 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0855 $X2=0.0270 $Y2=0.0360
r24 17 31 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0855 $X2=0.0270 $Y2=0.1350
r25 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2125 $Y2=0.0360
r26 27 28 11.7761 $w=1.3e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2125 $Y2=0.0360
r27 26 27 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r28 18 26 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r29 18 20 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r30 1 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r31 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r32 1 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r33 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r34 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AND3x4_ASAP7_75t_R%NET83 VSS 15 16 17 18 82 84 86 97 100 4 3 1 29 25
+ 24 20 26 6 19 21 5 28 22 30 23 31 27
c1 1 VSS 0.0170107f
c2 3 VSS 0.00802277f
c3 4 VSS 0.00828036f
c4 5 VSS 0.00447225f
c5 6 VSS 0.00807614f
c6 15 VSS 0.0808511f
c7 16 VSS 0.0800688f
c8 17 VSS 0.0803702f
c9 18 VSS 0.080593f
c10 19 VSS 0.00529687f
c11 20 VSS 0.00660712f
c12 21 VSS 0.00732871f
c13 22 VSS 0.00669804f
c14 23 VSS 0.00159976f
c15 24 VSS 0.00536272f
c16 25 VSS 0.00368972f
c17 26 VSS 0.0459915f
c18 27 VSS 0.00958939f
c19 28 VSS 0.0125123f
c20 29 VSS 0.000259642f
c21 30 VSS 0.00279263f
c22 31 VSS 0.00419696f
c23 32 VSS 0.00432081f
r1 100 99 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r2 5 99 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r3 96 5 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6380 $Y=0.0675 $X2=0.6500 $Y2=0.0675
r4 19 96 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6380 $Y2=0.0675
r5 97 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
r6 5 94 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r7 94 95 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.6480
+ $Y=0.0360 $X2=0.6790 $Y2=0.0360
r8 27 31 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7145
+ $Y=0.0360 $X2=0.7370 $Y2=0.0360
r9 27 95 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7145
+ $Y=0.0360 $X2=0.6790 $Y2=0.0360
r10 31 92 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.0360 $X2=0.7370 $Y2=0.0540
r11 91 92 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.0720 $X2=0.7370 $Y2=0.0540
r12 90 91 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.0900 $X2=0.7370 $Y2=0.0720
r13 89 90 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.1080 $X2=0.7370 $Y2=0.0900
r14 88 89 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.1530 $X2=0.7370 $Y2=0.1080
r15 87 88 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.1980 $X2=0.7370 $Y2=0.1530
r16 28 32 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.2160 $X2=0.7370 $Y2=0.2340
r17 28 87 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.2160 $X2=0.7370 $Y2=0.1980
r18 86 85 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r19 22 85 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6500 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r20 84 83 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r21 21 83 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r22 20 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r23 82 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r24 32 80 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.7370
+ $Y=0.2340 $X2=0.7145 $Y2=0.2340
r25 6 77 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6440 $Y2=0.2340
r26 4 72 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r27 3 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r28 79 80 8.27824 $w=1.3e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6790
+ $Y=0.2340 $X2=0.7145 $Y2=0.2340
r29 78 79 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6530
+ $Y=0.2340 $X2=0.6790 $Y2=0.2340
r30 77 78 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.6440
+ $Y=0.2340 $X2=0.6530 $Y2=0.2340
r31 76 77 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6255
+ $Y=0.2340 $X2=0.6440 $Y2=0.2340
r32 75 76 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5765
+ $Y=0.2340 $X2=0.6255 $Y2=0.2340
r33 74 75 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5225
+ $Y=0.2340 $X2=0.5765 $Y2=0.2340
r34 73 74 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.2340 $X2=0.5225 $Y2=0.2340
r35 72 73 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r36 71 72 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4745
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r37 70 71 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4745 $Y2=0.2340
r38 69 70 15.1573 $w=1.3e-08 $l=6.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r39 68 69 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r40 67 68 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r41 66 67 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r42 26 30 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.2690 $Y2=0.2340
r43 26 66 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2940
+ $Y=0.2340 $X2=0.3125 $Y2=0.2340
r44 30 65 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2690
+ $Y=0.2340 $X2=0.2690 $Y2=0.2160
r45 64 65 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2690
+ $Y=0.2035 $X2=0.2690 $Y2=0.2160
r46 25 29 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2690 $Y=0.1720 $X2=0.2690 $Y2=0.1350
r47 25 64 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2690
+ $Y=0.1720 $X2=0.2690 $Y2=0.2035
r48 24 29 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2690 $Y=0.0980 $X2=0.2690 $Y2=0.1350
r49 29 60 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2690 $Y=0.1350 $X2=0.2560 $Y2=0.1350
r50 59 60 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2560 $Y2=0.1350
r51 58 59 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r52 23 58 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2240
+ $Y=0.1350 $X2=0.2320 $Y2=0.1350
r53 18 52 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r54 17 45 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r55 16 39 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r56 52 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r57 51 52 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r58 49 51 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2335 $Y2=0.1350
r59 48 49 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r60 46 48 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2160 $Y2=0.1350
r61 45 46 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r62 43 45 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r63 42 43 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r64 40 42 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r65 39 40 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r66 37 39 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r67 36 37 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r68 35 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r69 15 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r70 1 34 3.20232 $w=2.13909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r71 1 35 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r72 15 34 0.905388 $w=2.07755e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0700 $Y2=0.1350
r73 15 35 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r74 6 22 1e-05
r75 4 21 1e-05
.ends

.subckt PM_AND3x4_ASAP7_75t_R%NET89 VSS 15 29 30 32 13 12 11 3 2 1 10
c1 1 VSS 0.00386872f
c2 2 VSS 0.00306194f
c3 3 VSS 0.00426211f
c4 10 VSS 0.00281613f
c5 11 VSS 0.0021011f
c6 12 VSS 0.00239345f
c7 13 VSS 0.00313339f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7000 $Y2=0.0675
r2 32 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r3 30 28 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r4 2 28 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5940 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5940 $Y2=0.0675
r6 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r7 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6960 $Y=0.0675
+ $X2=0.6920 $Y2=0.0720
r8 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0720
r9 25 26 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6660
+ $Y=0.0720 $X2=0.6920 $Y2=0.0720
r10 24 25 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6415
+ $Y=0.0720 $X2=0.6660 $Y2=0.0720
r11 23 24 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6230
+ $Y=0.0720 $X2=0.6415 $Y2=0.0720
r12 22 23 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6075
+ $Y=0.0720 $X2=0.6230 $Y2=0.0720
r13 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5940
+ $Y=0.0720 $X2=0.6075 $Y2=0.0720
r14 20 21 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5695
+ $Y=0.0720 $X2=0.5940 $Y2=0.0720
r15 19 20 5.13017 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.5475
+ $Y=0.0720 $X2=0.5695 $Y2=0.0720
r16 18 19 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5225
+ $Y=0.0720 $X2=0.5475 $Y2=0.0720
r17 17 18 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.0720 $X2=0.5225 $Y2=0.0720
r18 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0720 $X2=0.4995 $Y2=0.0720
r19 13 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4745
+ $Y=0.0720 $X2=0.4860 $Y2=0.0720
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0720
r21 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r22 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4880 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r23 1 10 1e-05
.ends


*
.SUBCKT AND3x4_ASAP7_75t_R VSS VDD C B A Y
*
* VSS VSS
* VDD VDD
* C C
* B B
* A A
* Y Y
*
*

MM7 N_MM7_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@4 N_MM7@4_d N_MM6@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@3 N_MM7@3_d N_MM6@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7@2 N_MM7@2_d N_MM6@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2@2 N_MM2@2_d N_MM2@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM4_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM3_g N_MM0@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@4 N_MM6@4_d N_MM6@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@3 N_MM6@3_d N_MM6@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND3x4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND3x4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND3x4_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND3x4_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM2@2_g 0.0016265f
cc_2 N_noxref_12_1 N_NET89_10 0.000589562f
x_PM_AND3x4_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AND3x4_ASAP7_75t_R%noxref_14
cc_3 N_noxref_14_1 N_MM4_g 0.00144531f
cc_4 N_noxref_14_1 N_NET89_10 0.0360711f
cc_5 N_noxref_14_1 N_noxref_12_1 0.00765663f
cc_6 N_noxref_14_1 N_noxref_13_1 0.000480998f
x_PM_AND3x4_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_AND3x4_ASAP7_75t_R%noxref_10
cc_7 N_noxref_10_1 N_MM7_g 0.00146202f
cc_8 N_noxref_10_1 N_Y_13 0.000837308f
x_PM_AND3x4_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_AND3x4_ASAP7_75t_R%noxref_11
cc_9 N_noxref_11_1 N_MM7_g 0.00146346f
cc_10 N_noxref_11_1 N_Y_15 0.000844065f
cc_11 N_noxref_11_1 N_noxref_10_1 0.00176462f
x_PM_AND3x4_ASAP7_75t_R%NET90 VSS N_MM2_d N_MM2@2_d N_MM1_s N_MM1@2_s N_NET90_9
+ N_NET90_7 N_NET90_1 N_NET90_2 N_NET90_8 PM_AND3x4_ASAP7_75t_R%NET90
cc_12 N_NET90_9 N_NET83_29 7.06091e-20
cc_13 N_NET90_9 N_NET83_26 0.000113443f
cc_14 N_NET90_9 N_NET83_4 0.000823693f
cc_15 N_NET90_9 N_NET83_24 0.00174337f
cc_16 N_NET90_7 N_C_1 0.00189608f
cc_17 N_NET90_1 N_C_5 0.0019258f
cc_18 N_NET90_1 N_MM2@2_g 0.00208031f
cc_19 N_NET90_7 N_MM5_g 0.0181291f
cc_20 N_NET90_7 N_MM2@2_g 0.0500279f
cc_21 N_NET90_2 N_MM1@2_g 0.00182661f
cc_22 N_NET90_8 N_B_1 0.0019965f
cc_23 N_NET90_8 N_MM4_g 0.018199f
cc_24 N_NET90_8 N_MM1@2_g 0.0492324f
x_PM_AND3x4_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AND3x4_ASAP7_75t_R%noxref_15
cc_25 N_noxref_15_1 N_NET83_4 0.000429877f
cc_26 N_noxref_15_1 N_NET83_21 0.0367152f
cc_27 N_noxref_15_1 N_MM4_g 0.00146142f
cc_28 N_noxref_15_1 N_noxref_13_1 0.00780807f
cc_29 N_noxref_15_1 N_noxref_14_1 0.00124108f
x_PM_AND3x4_ASAP7_75t_R%B VSS B N_MM4_g N_MM1@2_g N_B_5 N_B_1 N_B_7 N_B_6
+ PM_AND3x4_ASAP7_75t_R%B
cc_30 N_MM4_g N_NET83_4 0.00222236f
cc_31 N_MM4_g N_NET83_6 0.000166381f
cc_32 N_MM4_g N_NET83_19 0.000367172f
cc_33 N_B_5 N_NET83_4 0.000944714f
cc_34 N_B_1 N_NET83_21 0.00104245f
cc_35 N_B_7 N_NET83_26 0.00553005f
cc_36 N_MM4_g N_NET83_21 0.0351155f
x_PM_AND3x4_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AND3x4_ASAP7_75t_R%noxref_13
cc_37 N_noxref_13_1 N_NET83_4 0.000188451f
cc_38 N_noxref_13_1 N_NET83_26 0.000226143f
cc_39 N_noxref_13_1 N_NET83_21 0.00123552f
cc_40 N_noxref_13_1 N_MM2@2_g 0.00918721f
cc_41 N_noxref_13_1 N_MM4_g 0.000274862f
cc_42 N_noxref_13_1 N_noxref_12_1 0.0013584f
x_PM_AND3x4_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AND3x4_ASAP7_75t_R%noxref_17
cc_43 N_noxref_17_1 N_NET83_28 0.000350228f
cc_44 N_noxref_17_1 N_NET83_22 0.000588607f
cc_45 N_noxref_17_1 N_MM3_g 0.00146363f
cc_46 N_noxref_17_1 N_NET89_12 0.000488143f
cc_47 N_noxref_17_1 N_noxref_16_1 0.00177219f
x_PM_AND3x4_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AND3x4_ASAP7_75t_R%noxref_16
cc_48 N_noxref_16_1 N_NET83_28 0.00034761f
cc_49 N_noxref_16_1 N_NET83_19 0.000569613f
cc_50 N_noxref_16_1 N_MM3_g 0.00145866f
cc_51 N_noxref_16_1 N_NET89_12 0.0360566f
x_PM_AND3x4_ASAP7_75t_R%C VSS C N_MM5_g N_MM2@2_g N_C_5 N_C_1
+ PM_AND3x4_ASAP7_75t_R%C
cc_52 N_MM2@2_g N_NET83_4 0.000134848f
cc_53 N_MM2@2_g N_NET83_3 0.0032652f
cc_54 N_MM2@2_g N_NET83_1 0.000419775f
cc_55 N_MM2@2_g N_NET83_29 0.000426107f
cc_56 N_MM2@2_g N_NET83_25 0.000728471f
cc_57 N_MM2@2_g N_NET83_24 0.000763814f
cc_58 N_MM5_g N_NET83_20 0.0328816f
cc_59 N_MM5_g N_MM6@2_g 0.00167274f
cc_60 N_C_5 N_NET83_26 0.00190374f
cc_61 N_C_1 N_NET83_20 0.00316255f
cc_62 N_C_5 N_NET83_3 0.00361851f
cc_63 N_MM2@2_g N_NET83_20 0.0414694f
x_PM_AND3x4_ASAP7_75t_R%A VSS A N_MM0_g N_MM3_g N_A_5 N_A_1 N_A_7 N_A_6
+ PM_AND3x4_ASAP7_75t_R%A
cc_64 N_MM3_g N_NET83_6 0.00347186f
cc_65 N_MM3_g N_NET83_5 0.00239391f
cc_66 N_MM3_g N_NET83_28 0.000823991f
cc_67 N_A_5 N_NET83_6 0.00109044f
cc_68 N_MM3_g N_NET83_22 0.0335869f
cc_69 N_A_1 N_NET83_22 0.00429278f
cc_70 N_A_7 N_NET83_26 0.00599488f
cc_71 N_MM0_g N_NET83_19 0.0384995f
cc_72 N_MM3_g N_NET83_19 0.0694216f
cc_73 N_A_1 N_B_1 0.00148184f
cc_74 N_MM0_g N_MM1@2_g 0.0127479f
x_PM_AND3x4_ASAP7_75t_R%Y VSS Y N_MM7_d N_MM7@4_d N_MM7@3_d N_MM7@2_d N_MM6_d
+ N_MM6@4_d N_MM6@3_d N_MM6@2_d N_Y_13 N_Y_4 N_Y_15 N_Y_16 N_Y_14 N_Y_19 N_Y_18
+ N_Y_2 N_Y_1 N_Y_3 PM_AND3x4_ASAP7_75t_R%Y
cc_75 N_Y_13 N_NET83_24 0.00023725f
cc_76 N_Y_13 N_NET83_30 0.000779091f
cc_77 N_Y_13 N_NET83_1 0.00107319f
cc_78 N_Y_4 N_NET83_23 0.000830318f
cc_79 N_Y_15 N_MM6@4_g 0.0306162f
cc_80 N_Y_16 N_MM6@2_g 0.030666f
cc_81 N_Y_14 N_MM6@2_g 0.0673577f
cc_82 N_Y_19 N_NET83_25 0.000954086f
cc_83 N_Y_18 N_NET83_24 0.00115171f
cc_84 N_Y_18 N_MM6@4_g 0.00116487f
cc_85 N_Y_19 N_MM6@4_g 0.0013555f
cc_86 N_Y_2 N_MM6@4_g 0.00183839f
cc_87 N_Y_1 N_MM6@4_g 0.00188446f
cc_88 N_Y_3 N_MM6@2_g 0.00218269f
cc_89 N_Y_4 N_MM6@2_g 0.0022152f
cc_90 N_Y_15 N_NET83_1 0.00951519f
cc_91 N_Y_13 N_MM7_g 0.0367558f
cc_92 N_Y_14 N_MM6@3_g 0.0368809f
cc_93 N_Y_13 N_MM6@4_g 0.0678003f
x_PM_AND3x4_ASAP7_75t_R%NET83 VSS N_MM7_g N_MM6@4_g N_MM6@3_g N_MM6@2_g N_MM5_d
+ N_MM4_d N_MM3_d N_MM0_d N_MM0@2_d N_NET83_4 N_NET83_3 N_NET83_1 N_NET83_29
+ N_NET83_25 N_NET83_24 N_NET83_20 N_NET83_26 N_NET83_6 N_NET83_19 N_NET83_21
+ N_NET83_5 N_NET83_28 N_NET83_22 N_NET83_30 N_NET83_23 N_NET83_31 N_NET83_27
+ PM_AND3x4_ASAP7_75t_R%NET83
x_PM_AND3x4_ASAP7_75t_R%NET89 VSS N_MM1_d N_MM1@2_d N_MM0_s N_MM0@2_s
+ N_NET89_13 N_NET89_12 N_NET89_11 N_NET89_3 N_NET89_2 N_NET89_1 N_NET89_10
+ PM_AND3x4_ASAP7_75t_R%NET89
cc_94 N_NET89_13 N_NET83_31 0.000179165f
cc_95 N_NET89_13 N_NET83_21 0.000397311f
cc_96 N_NET89_13 N_NET83_4 0.000188494f
cc_97 N_NET89_13 N_NET83_26 0.00023289f
cc_98 N_NET89_13 N_NET83_5 0.00116764f
cc_99 N_NET89_12 N_NET83_19 0.000339769f
cc_100 N_NET89_11 N_NET83_19 0.000564242f
cc_101 N_NET89_3 N_NET83_27 0.000982451f
cc_102 N_NET89_2 N_NET83_5 0.00127389f
cc_103 N_NET89_3 N_NET83_19 0.00139756f
cc_104 N_NET89_3 N_NET83_28 0.00207935f
cc_105 N_NET89_3 N_NET83_5 0.00816414f
cc_106 N_NET89_13 N_NET83_27 0.00885661f
cc_107 N_NET89_2 N_MM1@2_g 0.000742648f
cc_108 N_NET89_1 N_MM4_g 0.00108055f
cc_109 N_NET89_11 N_B_1 0.00178995f
cc_110 N_NET89_13 N_B_6 0.00499245f
cc_111 N_NET89_11 N_MM1@2_g 0.0333611f
cc_112 N_NET89_10 N_MM4_g 0.0356502f
cc_113 N_NET89_2 N_MM3_g 0.00144186f
cc_114 N_NET89_3 N_MM3_g 0.00163009f
cc_115 N_NET89_3 N_A_1 0.00187337f
cc_116 N_NET89_13 N_A_6 0.00520691f
cc_117 N_NET89_11 N_MM0_g 0.0333388f
cc_118 N_NET89_12 N_MM3_g 0.0350133f
cc_119 N_NET89_1 N_NET90_9 0.000601234f
cc_120 N_NET89_13 N_NET90_2 0.00074454f
cc_121 N_NET89_11 N_NET90_8 0.00111907f
cc_122 N_NET89_1 N_NET90_2 0.00178534f
cc_123 N_NET89_2 N_NET90_2 0.00432272f
cc_124 N_NET89_13 N_NET90_9 0.0104011f
*END of AND3x4_ASAP7_75t_R.pxi
.ENDS
** Design:	AND4x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND4x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND4x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND4x1_ASAP7_75t_R%PD1 VSS 2 3 1
c1 1 VSS 0.000925075f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND4x1_ASAP7_75t_R%PD3 VSS 2 3 1
c1 1 VSS 0.000920533f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AND4x1_ASAP7_75t_R%PD2 VSS 2 3 1
c1 1 VSS 0.000914502f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AND4x1_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00522715f
c2 3 VSS 0.0457922f
c3 4 VSS 0.00705024f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_AND4x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0052678f
.ends

.subckt PM_AND4x1_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.0061646f
c2 3 VSS 0.0465571f
c3 4 VSS 0.0078896f
r1 8 4 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0800
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AND4x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0419661f
.ends

.subckt PM_AND4x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00464484f
.ends

.subckt PM_AND4x1_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00669732f
c2 3 VSS 0.045694f
c3 4 VSS 0.00471126f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_AND4x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00474198f
.ends

.subckt PM_AND4x1_ASAP7_75t_R%D VSS 10 3 4 1
c1 1 VSS 0.0065813f
c2 3 VSS 0.0835778f
c3 4 VSS 0.00930447f
r1 10 9 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1230
r2 4 9 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0825 $X2=0.2430 $Y2=0.1230
r3 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AND4x1_ASAP7_75t_R%Y VSS 18 14 27 7 1 2 8 9 10
c1 1 VSS 0.00959422f
c2 2 VSS 0.00803949f
c3 7 VSS 0.00379896f
c4 8 VSS 0.00373765f
c5 9 VSS 0.00419578f
c6 10 VSS 0.00381753f
c7 11 VSS 0.00656688f
c8 12 VSS 0.00290252f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r4 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r5 9 22 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r6 12 21 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3510 $Y2=0.2160
r7 12 23 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3375 $Y2=0.2340
r8 20 21 12.2425 $w=1.3e-08 $l=5.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1635 $X2=0.3510 $Y2=0.2160
r9 19 20 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1175 $X2=0.3510 $Y2=0.1635
r10 18 19 0.699569 $w=1.3e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1145 $X2=0.3510 $Y2=0.1175
r11 18 10 8.16164 $w=1.3e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1145 $X2=0.3510 $Y2=0.0795
r12 10 17 8.96345 $w=1.40345e-08 $l=4.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0795 $X2=0.3510 $Y2=0.0360
r13 16 17 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3375 $Y=0.0360 $X2=0.3510 $Y2=0.0360
r14 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r15 11 15 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r16 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r17 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r18 14 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
.ends

.subckt PM_AND4x1_ASAP7_75t_R%NET12 VSS 12 48 49 52 53 60 14 17 3 18 4 16 13 5
+ 24 15 20 1 21 26
c1 1 VSS 0.00329982f
c2 3 VSS 0.00595935f
c3 4 VSS 0.00995937f
c4 5 VSS 0.00996896f
c5 12 VSS 0.0800313f
c6 13 VSS 0.00319469f
c7 14 VSS 0.00491106f
c8 15 VSS 0.00492937f
c9 16 VSS 0.00538492f
c10 17 VSS 0.00495487f
c11 18 VSS 0.0183506f
c12 19 VSS 0.00060809f
c13 20 VSS 0.00137687f
c14 21 VSS 0.00127697f
c15 22 VSS 0.00290233f
c16 23 VSS 0.00343302f
c17 24 VSS 0.000509288f
c18 25 VSS 0.0027556f
c19 26 VSS 0.000595237f
r1 60 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r2 13 59 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r3 3 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r4 17 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r5 17 22 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r6 22 55 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r7 54 55 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.0575
r8 16 23 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2125 $X2=0.0270 $Y2=0.2340
r9 16 54 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2125 $X2=0.0270 $Y2=0.1350
r10 53 51 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r11 4 51 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r12 14 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r13 52 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r14 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r15 5 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r16 15 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r17 48 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r18 23 45 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0540 $Y2=0.2340
r19 4 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r20 5 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r21 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r22 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r23 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r24 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r25 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r26 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r27 38 39 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r28 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r29 18 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r30 18 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r31 25 37 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2340 $X2=0.2295 $Y2=0.2340
r32 19 35 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.2160 $X2=0.2430 $Y2=0.2035
r33 19 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2160 $X2=0.2430 $Y2=0.2340
r34 24 35 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1945 $X2=0.2430 $Y2=0.2035
r35 20 26 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r36 20 35 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1980 $X2=0.2430 $Y2=0.2035
r37 26 34 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1765
r38 33 34 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1540 $X2=0.2970 $Y2=0.1765
r39 32 33 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1540
r40 21 32 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1230 $X2=0.2970 $Y2=0.1350
r41 29 31 2.51167 $w=1.2975e-08 $l=2e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3085 $Y2=0.1350
r42 28 29 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r43 28 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r44 1 28 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r45 1 30 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r46 12 28 3.79335 $w=1.28e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r47 12 30 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r48 12 31 2.63307 $w=1.98865e-07 $l=1.15e-08 $layer=LIG $thickness=5.49565e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3085 $Y2=0.1350
r49 3 13 1e-05
.ends


*
.SUBCKT AND4x1_ASAP7_75t_R VSS VDD A B C D Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND4x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND4x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND4x1_ASAP7_75t_R%PD1 VSS N_MM0_s N_MM4_d N_PD1_1
+ PM_AND4x1_ASAP7_75t_R%PD1
cc_1 N_PD1_1 N_MM0_g 0.0172412f
cc_2 N_PD1_1 N_MM4_g 0.0172162f
x_PM_AND4x1_ASAP7_75t_R%PD3 VSS N_MM3_s N_MM5_d N_PD3_1
+ PM_AND4x1_ASAP7_75t_R%PD3
cc_3 N_PD3_1 N_MM3_g 0.0172996f
cc_4 N_PD3_1 N_MM5_g 0.0171839f
x_PM_AND4x1_ASAP7_75t_R%PD2 VSS N_MM4_s N_MM3_d N_PD2_1
+ PM_AND4x1_ASAP7_75t_R%PD2
cc_5 N_PD2_1 N_MM4_g 0.017382f
cc_6 N_PD2_1 N_MM3_g 0.0173278f
x_PM_AND4x1_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4 PM_AND4x1_ASAP7_75t_R%B
cc_7 N_B_1 N_A_1 0.00110928f
cc_8 N_MM4_g N_MM0_g 0.00515308f
cc_9 N_B_4 N_A_4 0.00657441f
x_PM_AND4x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND4x1_ASAP7_75t_R%noxref_12
cc_10 N_noxref_12_1 N_MM0_g 0.00145864f
cc_11 N_noxref_12_1 N_NET12_13 0.0379351f
x_PM_AND4x1_ASAP7_75t_R%C VSS C N_MM3_g N_C_1 N_C_4 PM_AND4x1_ASAP7_75t_R%C
cc_12 N_C_1 N_B_1 0.00113283f
cc_13 N_MM3_g N_MM4_g 0.00543369f
cc_14 N_C_4 N_B_4 0.00758745f
x_PM_AND4x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AND4x1_ASAP7_75t_R%noxref_13
cc_15 N_noxref_13_1 N_MM0_g 0.00145753f
cc_16 N_noxref_13_1 N_NET12_14 0.00131198f
cc_17 N_noxref_13_1 N_noxref_12_1 0.00178178f
x_PM_AND4x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AND4x1_ASAP7_75t_R%noxref_14
cc_18 N_noxref_14_1 N_MM9_g 0.00144579f
cc_19 N_noxref_14_1 N_Y_7 0.0385472f
x_PM_AND4x1_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_AND4x1_ASAP7_75t_R%A
x_PM_AND4x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AND4x1_ASAP7_75t_R%noxref_15
cc_20 N_noxref_15_1 N_MM9_g 0.00145848f
cc_21 N_noxref_15_1 N_Y_8 0.0384745f
cc_22 N_noxref_15_1 N_noxref_14_1 0.00177713f
x_PM_AND4x1_ASAP7_75t_R%D VSS D N_MM5_g N_D_4 N_D_1 PM_AND4x1_ASAP7_75t_R%D
cc_23 N_D_4 N_C_1 0.0010665f
cc_24 N_MM5_g N_MM3_g 0.0052216f
cc_25 N_D_4 N_C_4 0.00663611f
x_PM_AND4x1_ASAP7_75t_R%Y VSS Y N_MM9_d N_MM8_d N_Y_7 N_Y_1 N_Y_2 N_Y_8 N_Y_9
+ N_Y_10 PM_AND4x1_ASAP7_75t_R%Y
cc_26 N_Y_7 N_NET12_20 0.000396133f
cc_27 N_Y_7 N_NET12_1 0.000875843f
cc_28 N_Y_1 N_MM9_g 0.00105713f
cc_29 N_Y_2 N_MM9_g 0.0013982f
cc_30 N_Y_8 N_NET12_1 0.00146438f
cc_31 N_Y_9 N_NET12_26 0.00281881f
cc_32 N_Y_10 N_NET12_21 0.00464729f
cc_33 N_Y_8 N_MM9_g 0.0152508f
cc_34 N_Y_7 N_MM9_g 0.0553098f
x_PM_AND4x1_ASAP7_75t_R%NET12 VSS N_MM9_g N_MM2_d N_MM1_d N_MM7_d N_MM6_d
+ N_MM0_d N_NET12_14 N_NET12_17 N_NET12_3 N_NET12_18 N_NET12_4 N_NET12_16
+ N_NET12_13 N_NET12_5 N_NET12_24 N_NET12_15 N_NET12_20 N_NET12_1 N_NET12_21
+ N_NET12_26 PM_AND4x1_ASAP7_75t_R%NET12
cc_35 N_NET12_14 N_MM0_g 0.0157258f
cc_36 N_NET12_17 N_A_4 0.000754788f
cc_37 N_NET12_3 N_A_1 0.000956366f
cc_38 N_NET12_18 N_A_4 0.00107914f
cc_39 N_NET12_4 N_MM0_g 0.00115268f
cc_40 N_NET12_14 N_A_1 0.00140676f
cc_41 N_NET12_3 N_MM0_g 0.00168229f
cc_42 N_NET12_16 N_A_4 0.00830603f
cc_43 N_NET12_13 N_MM0_g 0.0547494f
cc_44 N_NET12_4 N_MM4_g 0.00150939f
cc_45 N_NET12_3 N_MM4_g 0.000330538f
cc_46 N_NET12_17 N_B_4 0.000387043f
cc_47 N_NET12_14 N_B_1 0.000637181f
cc_48 N_NET12_18 N_B_4 0.00115498f
cc_49 N_NET12_4 N_B_4 0.00248543f
cc_50 N_NET12_14 N_MM4_g 0.0357059f
cc_51 N_NET12_5 N_MM3_g 0.00145738f
cc_52 N_NET12_24 N_MM3_g 0.000366714f
cc_53 N_NET12_15 N_C_1 0.000688325f
cc_54 N_NET12_18 N_C_4 0.00109152f
cc_55 N_NET12_5 N_C_4 0.00245637f
cc_56 N_NET12_15 N_MM3_g 0.0354694f
cc_57 N_NET12_20 N_MM5_g 0.000381333f
cc_58 N_NET12_1 N_MM5_g 0.000445871f
cc_59 N_NET12_24 N_MM5_g 0.000526905f
cc_60 N_NET12_5 N_D_1 0.000663151f
cc_61 N_NET12_5 N_MM5_g 0.000950586f
cc_62 N_NET12_15 N_D_1 0.00102869f
cc_63 N_MM9_g N_MM5_g 0.00165279f
cc_64 N_NET12_21 N_D_4 0.00353533f
cc_65 N_NET12_15 N_MM5_g 0.0368215f
*END of AND4x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AND4x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND4x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND4x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND4x2_ASAP7_75t_R%NET17 VSS 2 3 1
c1 1 VSS 0.000926497f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_AND4x2_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000890704f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AND4x2_ASAP7_75t_R%NET15 VSS 2 3 1
c1 1 VSS 0.000938007f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AND4x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.042342f
.ends

.subckt PM_AND4x2_ASAP7_75t_R%D VSS 10 3 4 1
c1 1 VSS 0.00695183f
c2 3 VSS 0.0836175f
c3 4 VSS 0.00946012f
r1 10 9 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1225
r2 4 9 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0820 $X2=0.1890 $Y2=0.1225
r3 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_AND4x2_ASAP7_75t_R%A VSS 8 3 4 1
c1 1 VSS 0.00677444f
c2 3 VSS 0.0455756f
c3 4 VSS 0.00492638f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_AND4x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0423423f
.ends

.subckt PM_AND4x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00524552f
.ends

.subckt PM_AND4x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0419692f
.ends

.subckt PM_AND4x2_ASAP7_75t_R%Y VSS 21 16 17 28 29 7 8 11 9 2 1
c1 1 VSS 0.0117694f
c2 2 VSS 0.0100962f
c3 7 VSS 0.00459925f
c4 8 VSS 0.00452882f
c5 9 VSS 0.00741152f
c6 10 VSS 0.00974925f
c7 11 VSS 0.00888606f
c8 12 VSS 0.00340376f
c9 13 VSS 0.00345469f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 11 13 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r7 11 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r8 13 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r9 22 23 10.785 $w=1.3e-08 $l=4.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1697 $X2=0.0270 $Y2=0.2160
r10 21 22 8.80291 $w=1.3e-08 $l=3.77e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1320 $X2=0.0270 $Y2=0.1697
r11 21 20 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1320 $X2=0.0270 $Y2=0.1252
r12 9 12 9.07762 $w=1.49174e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0820 $X2=0.0270 $Y2=0.0360
r13 9 20 10.0855 $w=1.3e-08 $l=4.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0820 $X2=0.0270 $Y2=0.1252
r14 12 18 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0675 $Y2=0.0360
r15 10 18 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r16 1 10 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r17 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r18 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r20 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AND4x2_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00568215f
c2 3 VSS 0.0459566f
c3 4 VSS 0.00747066f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_AND4x2_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00549114f
c2 3 VSS 0.0463445f
c3 4 VSS 0.00786525f
r1 8 4 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0800
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_AND4x2_ASAP7_75t_R%NET33 VSS 12 13 56 57 60 61 68 20 23 1 3 17 15 21
+ 4 5 16 25 14 24 22 18
c1 1 VSS 0.0074137f
c2 3 VSS 0.00986895f
c3 4 VSS 0.00997465f
c4 5 VSS 0.0065478f
c5 12 VSS 0.081167f
c6 13 VSS 0.0808642f
c7 14 VSS 0.00493758f
c8 15 VSS 0.00653216f
c9 16 VSS 0.00654241f
c10 17 VSS 0.00219821f
c11 18 VSS 0.00118241f
c12 19 VSS 0.000692046f
c13 20 VSS 0.0226968f
c14 21 VSS 0.00903316f
c15 22 VSS 0.000464578f
c16 23 VSS 0.000913725f
c17 24 VSS 0.00276825f
c18 25 VSS 0.00693629f
c19 26 VSS 0.00395896f
r1 14 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3760 $Y2=0.0675
r2 68 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r3 5 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r4 65 66 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r5 25 63 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.4050 $Y2=0.0575
r6 25 66 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3915 $Y2=0.0360
r7 62 63 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.0575
r8 21 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2125 $X2=0.4050 $Y2=0.2340
r9 21 62 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2125 $X2=0.4050 $Y2=0.1350
r10 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r11 4 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r12 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r13 60 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r14 57 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r15 3 55 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r16 15 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r17 56 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r18 26 53 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.3800 $Y2=0.2340
r19 4 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r20 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r21 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.2340 $X2=0.3800 $Y2=0.2340
r22 51 52 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.2340 $X2=0.3620 $Y2=0.2340
r23 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.2340 $X2=0.3510 $Y2=0.2340
r24 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r25 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r26 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2340 $X2=0.3105 $Y2=0.2340
r27 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2970 $Y2=0.2340
r28 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r29 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r30 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2295 $Y2=0.2340
r31 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r32 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.2025 $Y2=0.2340
r33 20 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1755 $Y=0.2340 $X2=0.1620 $Y2=0.2340
r34 20 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r35 19 40 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.2160 $X2=0.1620 $Y2=0.2035
r36 19 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2160 $X2=0.1620 $Y2=0.2340
r37 23 40 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1945 $X2=0.1620 $Y2=0.2035
r38 39 40 3.9716 $w=1.39211e-08 $l=2.51098e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1375 $Y=0.1980 $X2=0.1620 $Y2=0.2035
r39 18 22 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1195 $Y=0.1980 $X2=0.1080 $Y2=0.1980
r40 18 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.1980 $X2=0.1375 $Y2=0.1980
r41 22 37 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1980 $X2=0.1080 $Y2=0.1765
r42 13 33 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r43 36 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1540 $X2=0.1080 $Y2=0.1765
r44 35 36 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1350 $X2=0.1080 $Y2=0.1540
r45 17 35 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1225 $X2=0.1080 $Y2=0.1350
r46 31 33 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r47 30 31 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r48 30 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1080 $Y=0.1350
+ $X2=0.1080 $Y2=0.1350
r49 29 30 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r50 12 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r51 1 28 4.63801 $w=1.7681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r52 1 29 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r53 12 28 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r54 12 29 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT AND4x2_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g N_MM8_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM4_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM5_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND4x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND4x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND4x2_ASAP7_75t_R%NET17 VSS N_MM7_d N_MM6_s N_NET17_1
+ PM_AND4x2_ASAP7_75t_R%NET17
cc_1 N_NET17_1 N_MM4_g 0.0172941f
cc_2 N_NET17_1 N_MM5_g 0.0171621f
x_PM_AND4x2_ASAP7_75t_R%NET16 VSS N_MM8_d N_MM7_s N_NET16_1
+ PM_AND4x2_ASAP7_75t_R%NET16
cc_3 N_NET16_1 N_MM8_g 0.0173911f
cc_4 N_NET16_1 N_MM4_g 0.0173438f
x_PM_AND4x2_ASAP7_75t_R%NET15 VSS N_MM9_d N_MM8_s N_NET15_1
+ PM_AND4x2_ASAP7_75t_R%NET15
cc_5 N_NET15_1 N_MM9_g 0.0172356f
cc_6 N_NET15_1 N_MM8_g 0.0172308f
x_PM_AND4x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_AND4x2_ASAP7_75t_R%noxref_12
cc_7 N_noxref_12_1 N_MM0_g 0.00147308f
cc_8 N_noxref_12_1 N_Y_7 0.000830204f
x_PM_AND4x2_ASAP7_75t_R%D VSS D N_MM9_g N_D_4 N_D_1 PM_AND4x2_ASAP7_75t_R%D
cc_9 N_MM9_g N_NET33_20 0.000217947f
cc_10 N_MM9_g N_NET33_23 0.000445898f
cc_11 N_MM9_g N_NET33_1 0.000537956f
cc_12 N_MM9_g N_NET33_3 0.00152674f
cc_13 N_D_4 N_NET33_17 0.000564826f
cc_14 N_D_1 N_NET33_15 0.00101098f
cc_15 N_MM9_g N_MM0@2_g 0.00165664f
cc_16 N_D_4 N_NET33_1 0.00170566f
cc_17 N_MM9_g N_NET33_15 0.036941f
x_PM_AND4x2_ASAP7_75t_R%A VSS A N_MM5_g N_A_4 N_A_1 PM_AND4x2_ASAP7_75t_R%A
cc_18 N_MM5_g N_NET33_16 0.0157014f
cc_19 N_A_4 N_NET33_25 0.000570539f
cc_20 N_A_1 N_NET33_5 0.000903332f
cc_21 N_A_4 N_NET33_20 0.0011516f
cc_22 N_MM5_g N_NET33_4 0.00121131f
cc_23 N_A_1 N_NET33_16 0.00145529f
cc_24 N_MM5_g N_NET33_5 0.00167152f
cc_25 N_A_4 N_NET33_21 0.00805763f
cc_26 N_MM5_g N_NET33_14 0.0547142f
cc_27 N_A_1 N_B_1 0.00118768f
cc_28 N_MM5_g N_MM4_g 0.00520938f
cc_29 N_A_4 N_B_4 0.00640562f
x_PM_AND4x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_AND4x2_ASAP7_75t_R%noxref_13
cc_30 N_noxref_13_1 N_MM0_g 0.00147501f
cc_31 N_noxref_13_1 N_Y_8 0.000834152f
cc_32 N_noxref_13_1 N_noxref_12_1 0.00177715f
x_PM_AND4x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AND4x2_ASAP7_75t_R%noxref_14
cc_33 N_noxref_14_1 N_NET33_5 0.000506524f
cc_34 N_noxref_14_1 N_NET33_14 0.0374608f
cc_35 N_noxref_14_1 N_MM5_g 0.00145668f
x_PM_AND4x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AND4x2_ASAP7_75t_R%noxref_15
cc_36 N_noxref_15_1 N_NET33_16 0.0013148f
cc_37 N_noxref_15_1 N_MM5_g 0.00145726f
cc_38 N_noxref_15_1 N_noxref_14_1 0.00177642f
x_PM_AND4x2_ASAP7_75t_R%Y VSS Y N_MM0_d N_MM0@2_d N_MM1_d N_MM1@2_d N_Y_7 N_Y_8
+ N_Y_11 N_Y_9 N_Y_2 N_Y_1 PM_AND4x2_ASAP7_75t_R%Y
cc_39 N_Y_7 N_NET33_17 0.000318771f
cc_40 N_Y_7 N_NET33_24 0.000343836f
cc_41 N_Y_7 N_NET33_22 0.000471081f
cc_42 N_Y_7 N_NET33_1 0.000865675f
cc_43 N_Y_8 N_MM0_g 0.0306345f
cc_44 N_Y_11 N_NET33_18 0.000956932f
cc_45 N_Y_9 N_NET33_1 0.00139688f
cc_46 N_Y_2 N_NET33_17 0.00183212f
cc_47 N_Y_1 N_MM0_g 0.00186432f
cc_48 N_Y_2 N_MM0_g 0.00248196f
cc_49 N_Y_11 N_NET33_22 0.00327101f
cc_50 N_Y_8 N_NET33_1 0.00426928f
cc_51 N_Y_7 N_MM0@2_g 0.0370928f
cc_52 N_Y_7 N_MM0_g 0.0683678f
x_PM_AND4x2_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4 PM_AND4x2_ASAP7_75t_R%B
cc_53 N_MM4_g N_NET33_21 0.000210741f
cc_54 N_MM4_g N_NET33_4 0.00149219f
cc_55 N_MM4_g N_NET33_5 0.000344731f
cc_56 N_B_1 N_NET33_16 0.000711123f
cc_57 N_B_4 N_NET33_20 0.0011926f
cc_58 N_B_4 N_NET33_4 0.00232326f
cc_59 N_MM4_g N_NET33_16 0.0356436f
cc_60 N_B_1 N_C_1 0.00128681f
cc_61 N_MM4_g N_MM8_g 0.00542776f
cc_62 N_B_4 N_C_4 0.00759022f
x_PM_AND4x2_ASAP7_75t_R%C VSS C N_MM8_g N_C_1 N_C_4 PM_AND4x2_ASAP7_75t_R%C
cc_63 N_MM8_g N_NET33_3 0.00149016f
cc_64 N_C_1 N_NET33_15 0.000551379f
cc_65 N_C_4 N_NET33_20 0.00128722f
cc_66 N_C_4 N_NET33_3 0.00217965f
cc_67 N_MM8_g N_NET33_15 0.0353397f
cc_68 N_C_1 N_D_4 0.00108091f
cc_69 N_MM8_g N_MM9_g 0.00522091f
cc_70 N_C_4 N_D_4 0.00676751f
x_PM_AND4x2_ASAP7_75t_R%NET33 VSS N_MM0_g N_MM0@2_g N_MM2_d N_MM3_d N_MM4_d
+ N_MM5_d N_MM6_d N_NET33_20 N_NET33_23 N_NET33_1 N_NET33_3 N_NET33_17
+ N_NET33_15 N_NET33_21 N_NET33_4 N_NET33_5 N_NET33_16 N_NET33_25 N_NET33_14
+ N_NET33_24 N_NET33_22 N_NET33_18 PM_AND4x2_ASAP7_75t_R%NET33
*END of AND4x2_ASAP7_75t_R.pxi
.ENDS
** Design:	AND5x1_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND5x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND5x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND5x1_ASAP7_75t_R%NET024 VSS 2 3 1
c1 1 VSS 0.00089714f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_AND5x1_ASAP7_75t_R%NET023 VSS 2 3 1
c1 1 VSS 0.000851318f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_AND5x1_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000860325f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_AND5x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000860487f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2700 $Y2=0.0675
.ends

.subckt PM_AND5x1_ASAP7_75t_R%B VSS 10 3 1 4
c1 1 VSS 0.00353131f
c2 3 VSS 0.0349253f
c3 4 VSS 0.00689588f
r1 10 9 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1340 $X2=0.1350 $Y2=0.0975
r2 4 9 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0575 $X2=0.1350 $Y2=0.0975
r3 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1345
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1340
+ $X2=0.1350 $Y2=0.1345
.ends

.subckt PM_AND5x1_ASAP7_75t_R%A VSS 8 3 1 4
c1 1 VSS 0.00472752f
c2 3 VSS 0.034431f
c3 4 VSS 0.00436195f
r1 8 4 8.51143 $w=1.3e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1340 $X2=0.0810 $Y2=0.0975
r2 3 1 3.49039 $w=1.235e-07 $l=1e-09 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1340
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1340
+ $X2=0.0810 $Y2=0.1340
.ends

.subckt PM_AND5x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00473774f
.ends

.subckt PM_AND5x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00480129f
.ends

.subckt PM_AND5x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.004408f
.ends

.subckt PM_AND5x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00458179f
.ends

.subckt PM_AND5x1_ASAP7_75t_R%E VSS 10 3 1 4
c1 1 VSS 0.0068927f
c2 3 VSS 0.0831891f
c3 4 VSS 0.00759844f
r1 10 9 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1340 $X2=0.2970 $Y2=0.1205
r2 4 9 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0805 $X2=0.2970 $Y2=0.1205
r3 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1345
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1340
+ $X2=0.2970 $Y2=0.1345
.ends

.subckt PM_AND5x1_ASAP7_75t_R%D VSS 8 3 1 4
c1 1 VSS 0.00420347f
c2 3 VSS 0.0355217f
c3 4 VSS 0.00766332f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1340 $X2=0.2430 $Y2=0.0795
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1345
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1340
+ $X2=0.2430 $Y2=0.1345
.ends

.subckt PM_AND5x1_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00374422f
c2 3 VSS 0.0350978f
c3 4 VSS 0.00681354f
r1 8 4 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1340 $X2=0.1890 $Y2=0.0795
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1345
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1340
+ $X2=0.1890 $Y2=0.1345
.ends

.subckt PM_AND5x1_ASAP7_75t_R%Y VSS 20 15 27 10 7 1 2 9 11 8
c1 1 VSS 0.00812816f
c2 2 VSS 0.00801046f
c3 7 VSS 0.00385536f
c4 8 VSS 0.00384419f
c5 9 VSS 0.00478699f
c6 10 VSS 0.00496925f
c7 11 VSS 0.00380717f
c8 12 VSS 0.0028477f
c9 13 VSS 0.00286929f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r4 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r5 9 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r6 13 22 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4050 $Y2=0.2160
r7 13 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.3915 $Y2=0.2340
r8 21 22 11.1348 $w=1.3e-08 $l=4.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1682 $X2=0.4050 $Y2=0.2160
r9 20 21 9.1527 $w=1.3e-08 $l=3.92e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1290 $X2=0.4050 $Y2=0.1682
r10 20 19 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1290 $X2=0.4050 $Y2=0.1222
r11 11 12 8.72783 $w=1.4982e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0805 $X2=0.4050 $Y2=0.0360
r12 11 19 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0805 $X2=0.4050 $Y2=0.1222
r13 12 17 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3915 $Y2=0.0360
r14 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r15 10 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r16 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r17 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3760 $Y2=0.0675
r18 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
.ends

.subckt PM_AND5x1_ASAP7_75t_R%NET011 VSS 15 54 55 58 59 63 68 25 4 3 21 16 17
+ 20 5 18 6 27 19 23 1 24 29
c1 1 VSS 0.00357793f
c2 3 VSS 0.00601675f
c3 4 VSS 0.00694027f
c4 5 VSS 0.00836223f
c5 6 VSS 0.0087625f
c6 15 VSS 0.0800278f
c7 16 VSS 0.00321015f
c8 17 VSS 0.00360804f
c9 18 VSS 0.00436272f
c10 19 VSS 0.00447261f
c11 20 VSS 0.00407353f
c12 21 VSS 0.0224968f
c13 22 VSS 0.00053735f
c14 23 VSS 0.0013644f
c15 24 VSS 0.00143734f
c16 25 VSS 0.00660076f
c17 26 VSS 0.00301037f
c18 27 VSS 0.000546338f
c19 28 VSS 0.00273513f
c20 29 VSS 0.000478736f
r1 68 67 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r2 16 67 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r3 3 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r4 64 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r5 25 61 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r6 25 64 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r7 63 62 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r8 17 62 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2160 $X2=0.0685 $Y2=0.2160
r9 60 61 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.0575
r10 20 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2125 $X2=0.0270 $Y2=0.2340
r11 20 60 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2125 $X2=0.0270 $Y2=0.1350
r12 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r13 5 57 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2160 $X2=0.1765 $Y2=0.2160
r14 18 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2160 $X2=0.1620 $Y2=0.2160
r15 58 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2160 $X2=0.1475 $Y2=0.2160
r16 54 53 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r17 6 53 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2160 $X2=0.2845 $Y2=0.2160
r18 19 6 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2160 $X2=0.2700 $Y2=0.2160
r19 55 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2160 $X2=0.2555 $Y2=0.2160
r20 4 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2160
+ $X2=0.0540 $Y2=0.2340
r21 26 49 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r22 5 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2160
+ $X2=0.1620 $Y2=0.2340
r23 6 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r24 50 51 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0665 $Y2=0.2340
r25 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r26 48 51 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0710
+ $Y=0.2340 $X2=0.0665 $Y2=0.2340
r27 47 48 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0710 $Y2=0.2340
r28 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r29 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r30 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r31 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r32 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r33 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1755 $Y2=0.2340
r34 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r35 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r36 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2835 $Y2=0.2340
r37 21 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r38 21 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r39 28 38 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2835 $Y2=0.2340
r40 22 36 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2160 $X2=0.2970 $Y2=0.2035
r41 22 28 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.2160 $X2=0.2970 $Y2=0.2340
r42 27 36 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1945 $X2=0.2970 $Y2=0.2035
r43 23 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.3510 $Y2=0.1980
r44 23 36 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.2970 $Y2=0.2035
r45 29 35 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1765
r46 34 35 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1535 $X2=0.3510 $Y2=0.1765
r47 33 34 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1340 $X2=0.3510 $Y2=0.1535
r48 24 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1205 $X2=0.3510 $Y2=0.1340
r49 15 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1345
r50 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1345
+ $X2=0.3510 $Y2=0.1340
r51 3 16 1e-05
r52 4 17 1e-05
.ends


*
.SUBCKT AND5x1_ASAP7_75t_R VSS VDD A B C D E Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* E E
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 N_MM2_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 N_MM7_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 N_MM8_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND5x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND5x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND5x1_ASAP7_75t_R%NET024 VSS N_MM0_s N_MM4_d N_NET024_1
+ PM_AND5x1_ASAP7_75t_R%NET024
cc_1 N_NET024_1 N_MM0_g 0.0174435f
cc_2 N_NET024_1 N_MM4_g 0.0174207f
x_PM_AND5x1_ASAP7_75t_R%NET023 VSS N_MM4_s N_MM3_d N_NET023_1
+ PM_AND5x1_ASAP7_75t_R%NET023
cc_3 N_NET023_1 N_MM4_g 0.0176216f
cc_4 N_NET023_1 N_MM3_g 0.0175335f
x_PM_AND5x1_ASAP7_75t_R%NET30 VSS N_MM3_s N_MM5_d N_NET30_1
+ PM_AND5x1_ASAP7_75t_R%NET30
cc_5 N_NET30_1 N_MM3_g 0.017636f
cc_6 N_NET30_1 N_MM5_g 0.0175099f
x_PM_AND5x1_ASAP7_75t_R%NET29 VSS N_MM5_s N_MM6_d N_NET29_1
+ PM_AND5x1_ASAP7_75t_R%NET29
cc_7 N_NET29_1 N_MM5_g 0.0175104f
cc_8 N_NET29_1 N_MM9_g 0.0173605f
x_PM_AND5x1_ASAP7_75t_R%B VSS B N_MM4_g N_B_1 N_B_4 PM_AND5x1_ASAP7_75t_R%B
cc_9 N_B_1 N_A_1 0.00143655f
cc_10 N_B_4 N_A_4 0.00555721f
cc_11 N_MM4_g N_MM0_g 0.00841497f
x_PM_AND5x1_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_AND5x1_ASAP7_75t_R%A
x_PM_AND5x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AND5x1_ASAP7_75t_R%noxref_16
cc_12 N_noxref_16_1 N_MM1_g 0.00145459f
cc_13 N_noxref_16_1 N_Y_7 0.0384575f
x_PM_AND5x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AND5x1_ASAP7_75t_R%noxref_14
cc_14 N_noxref_14_1 N_MM0_g 0.00160349f
cc_15 N_noxref_14_1 N_NET011_3 0.000509405f
cc_16 N_noxref_14_1 N_NET011_16 0.0376819f
x_PM_AND5x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AND5x1_ASAP7_75t_R%noxref_15
cc_17 N_noxref_15_1 N_MM0_g 0.00348451f
cc_18 N_noxref_15_1 N_NET011_4 0.000505215f
cc_19 N_noxref_15_1 N_NET011_17 0.0283488f
cc_20 N_noxref_15_1 N_noxref_14_1 0.00189799f
x_PM_AND5x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AND5x1_ASAP7_75t_R%noxref_17
cc_21 N_noxref_17_1 N_MM1_g 0.00145827f
cc_22 N_noxref_17_1 N_Y_8 0.0385852f
cc_23 N_noxref_17_1 N_noxref_16_1 0.00177677f
x_PM_AND5x1_ASAP7_75t_R%E VSS E N_MM9_g N_E_1 N_E_4 PM_AND5x1_ASAP7_75t_R%E
cc_24 N_E_1 N_D_1 0.00165692f
cc_25 N_E_4 N_D_4 0.00555868f
cc_26 N_MM9_g N_MM5_g 0.0083989f
x_PM_AND5x1_ASAP7_75t_R%D VSS D N_MM5_g N_D_1 N_D_4 PM_AND5x1_ASAP7_75t_R%D
cc_27 N_D_1 N_C_1 0.0016259f
cc_28 N_D_4 N_C_4 0.0065339f
cc_29 N_MM5_g N_MM3_g 0.00870579f
x_PM_AND5x1_ASAP7_75t_R%C VSS C N_MM3_g N_C_1 N_C_4 PM_AND5x1_ASAP7_75t_R%C
cc_30 N_C_1 N_B_1 0.0014966f
cc_31 N_C_4 N_B_4 0.00627502f
cc_32 N_MM3_g N_MM4_g 0.00866703f
x_PM_AND5x1_ASAP7_75t_R%Y VSS Y N_MM11_d N_MM1_d N_Y_10 N_Y_7 N_Y_1 N_Y_2 N_Y_9
+ N_Y_11 N_Y_8 PM_AND5x1_ASAP7_75t_R%Y
cc_33 N_Y_10 N_E_4 0.00196531f
cc_34 N_Y_7 N_NET011_29 0.000180589f
cc_35 N_Y_7 N_NET011_23 0.000456263f
cc_36 N_Y_1 N_NET011_1 0.000855138f
cc_37 N_Y_1 N_MM1_g 0.00104833f
cc_38 N_Y_2 N_MM1_g 0.00139631f
cc_39 N_Y_7 N_NET011_1 0.0015291f
cc_40 N_Y_9 N_NET011_29 0.00241709f
cc_41 N_Y_11 N_NET011_24 0.00467804f
cc_42 N_Y_8 N_MM1_g 0.0153825f
cc_43 N_Y_7 N_MM1_g 0.0549759f
x_PM_AND5x1_ASAP7_75t_R%NET011 VSS N_MM1_g N_MM9_d N_MM8_d N_MM2_d N_MM7_d
+ N_MM10_d N_MM0_d N_NET011_25 N_NET011_4 N_NET011_3 N_NET011_21 N_NET011_16
+ N_NET011_17 N_NET011_20 N_NET011_5 N_NET011_18 N_NET011_6 N_NET011_27
+ N_NET011_19 N_NET011_23 N_NET011_1 N_NET011_24 N_NET011_29
+ PM_AND5x1_ASAP7_75t_R%NET011
cc_44 N_NET011_25 N_A_4 0.000581549f
cc_45 N_NET011_4 N_MM0_g 0.000711449f
cc_46 N_NET011_3 N_A_1 0.000750565f
cc_47 N_NET011_21 N_A_4 0.00120676f
cc_48 N_NET011_16 N_A_1 0.00135405f
cc_49 N_NET011_3 N_MM0_g 0.00176143f
cc_50 N_NET011_17 N_MM0_g 0.0108577f
cc_51 N_NET011_20 N_A_4 0.00825983f
cc_52 N_NET011_16 N_MM0_g 0.0500341f
cc_53 N_NET011_25 N_MM4_g 0.000197444f
cc_54 N_NET011_20 N_MM4_g 0.000211253f
cc_55 N_NET011_3 N_MM4_g 0.000344075f
cc_56 N_NET011_5 N_MM4_g 0.000703504f
cc_57 N_NET011_21 N_B_4 0.00124854f
cc_58 N_NET011_3 N_B_4 0.00222208f
cc_59 N_NET011_18 N_MM4_g 0.0262197f
cc_60 N_NET011_5 N_MM3_g 0.000704974f
cc_61 N_NET011_21 N_C_4 0.00128757f
cc_62 N_NET011_5 N_C_4 0.00169215f
cc_63 N_NET011_18 N_MM3_g 0.0258086f
cc_64 N_NET011_6 N_MM5_g 0.000695822f
cc_65 N_NET011_21 N_D_4 0.00120719f
cc_66 N_NET011_27 N_D_4 0.00252639f
cc_67 N_NET011_19 N_MM5_g 0.0261236f
cc_68 N_NET011_23 N_MM9_g 0.000385408f
cc_69 N_NET011_6 N_MM9_g 0.000407182f
cc_70 N_NET011_27 N_MM9_g 0.000535038f
cc_71 N_NET011_1 N_E_1 0.00212866f
cc_72 N_NET011_24 N_E_4 0.00363574f
cc_73 N_NET011_19 N_MM9_g 0.0109303f
cc_74 N_MM1_g N_MM9_g 0.017482f
*END of AND5x1_ASAP7_75t_R.pxi
.ENDS
** Design:	AND5x2_ASAP7_75t_R
* Created:	"Thu Aug 16 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "AND5x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "AND5x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_AND5x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0420011f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00596513f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00736251f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0424189f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%NET33 VSS 11 14 23 26 1 7 2 8 9
c1 1 VSS 0.0106003f
c2 2 VSS 0.00485738f
c3 7 VSS 0.00476827f
c4 8 VSS 0.0023335f
c5 9 VSS 0.0267076f
r1 26 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r2 24 25 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3340 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r3 2 24 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3220 $Y=0.0675 $X2=0.3340 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r5 23 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r6 2 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r7 19 20 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r8 18 19 19.4713 $w=1.3e-08 $l=8.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2020
+ $Y=0.0360 $X2=0.2855 $Y2=0.0360
r9 17 18 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1325
+ $Y=0.0360 $X2=0.2020 $Y2=0.0360
r10 16 17 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1325 $Y2=0.0360
r11 15 16 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r12 9 15 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.0970 $Y2=0.0360
r13 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r14 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r15 1 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1100 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r16 10 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0980 $Y=0.0675 $X2=0.1100 $Y2=0.0675
r17 7 10 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.0980 $Y2=0.0675
r18 11 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_22 VSS 1
c1 1 VSS 0.00696415f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.00652144f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_23 VSS 1
c1 1 VSS 0.00577373f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%Y VSS 22 16 17 28 29 7 2 8 11 1
c1 1 VSS 0.0106236f
c2 2 VSS 0.0105881f
c3 7 VSS 0.00452723f
c4 8 VSS 0.00457202f
c5 9 VSS 0.00959032f
c6 10 VSS 0.00893315f
c7 11 VSS 0.0078618f
c8 12 VSS 0.00342062f
c9 13 VSS 0.00347006f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.2025 $X2=0.9865 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9720 $Y=0.2025 $X2=0.9865 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.2025 $X2=0.9720 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.2025 $X2=0.9575 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9720 $Y=0.2025
+ $X2=0.9720 $Y2=0.2340
r6 24 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.2340 $X2=1.0125 $Y2=0.2340
r7 10 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9605
+ $Y=0.2340 $X2=0.9720 $Y2=0.2340
r8 13 23 9.4274 $w=1.48568e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0530 $Y2=0.1865
r9 13 25 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.2340 $X2=1.0125 $Y2=0.2340
r10 22 23 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1475 $X2=1.0530 $Y2=0.1865
r11 22 21 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1475 $X2=1.0530 $Y2=0.1455
r12 20 21 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.1350 $X2=1.0530 $Y2=0.1455
r13 11 12 9.89378 $w=1.47818e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0855 $X2=1.0530 $Y2=0.0360
r14 11 20 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.0530
+ $Y=0.0855 $X2=1.0530 $Y2=0.1350
r15 12 19 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.0530 $Y=0.0360 $X2=1.0125 $Y2=0.0360
r16 18 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.9720
+ $Y=0.0360 $X2=1.0125 $Y2=0.0360
r17 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.9605
+ $Y=0.0360 $X2=0.9720 $Y2=0.0360
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.9720 $Y=0.0675
+ $X2=0.9720 $Y2=0.0360
r19 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9890 $Y=0.0675 $X2=0.9865 $Y2=0.0675
r20 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9720 $Y=0.0675 $X2=0.9865 $Y2=0.0675
r21 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.9575 $Y=0.0675 $X2=0.9720 $Y2=0.0675
r22 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.9550 $Y=0.0675 $X2=0.9575 $Y2=0.0675
.ends

.subckt PM_AND5x2_ASAP7_75t_R%A VSS 18 3 4 5 1 7 6
c1 1 VSS 0.00909578f
c2 3 VSS 0.00907823f
c3 4 VSS 0.0462349f
c4 5 VSS 0.00445088f
c5 6 VSS 0.00385169f
c6 7 VSS 0.00428028f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1980 $X2=0.7290 $Y2=0.1665
r2 18 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1665
r3 18 5 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1215
r4 5 6 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.7290 $Y=0.1215 $X2=0.7290 $Y2=0.1080
r5 3 14 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7290 $Y2=0.1350
r6 14 15 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.7290
+ $Y=0.1350 $X2=0.7385 $Y2=0.1350
r7 18 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.7290 $Y=0.1350
+ $X2=0.7290 $Y2=0.1350
r8 11 15 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.7415 $Y=0.1350 $X2=0.7385 $Y2=0.1350
r9 10 11 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7560 $Y=0.1350 $X2=0.7415 $Y2=0.1350
r10 9 10 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7705 $Y=0.1350 $X2=0.7560 $Y2=0.1350
r11 4 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.7830
+ $Y=0.1350 $X2=0.7830 $Y2=0.1350
r12 1 9 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7705 $Y2=0.1350
r13 1 17 3.67391 $w=1.9681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7935 $Y2=0.1350
r14 4 9 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7705 $Y2=0.1350
r15 4 17 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.7830 $Y=0.1350 $X2=0.7935 $Y2=0.1350
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0422377f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%E VSS 18 3 4 1
c1 1 VSS 0.00995631f
c2 3 VSS 0.0824888f
c3 4 VSS 0.080903f
c4 5 VSS 0.0140801f
c5 6 VSS 0.0137791f
c6 7 VSS 0.00489748f
c7 8 VSS 0.0026023f
r1 6 8 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r2 5 8 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1215 $X2=0.0270 $Y2=0.1350
r3 4 16 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r4 18 7 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0540 $Y2=0.1350
r5 7 8 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.1350 $X2=0.0270 $Y2=0.1350
r6 14 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r7 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r8 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r9 10 12 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r10 9 10 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r11 18 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r12 1 9 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r13 1 11 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r14 3 9 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r15 3 11 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r16 3 12 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0055667f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_24 VSS 1
c1 1 VSS 0.00678137f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%D VSS 5 3 4 1 7 6
c1 1 VSS 0.0121213f
c2 3 VSS 0.0460548f
c3 4 VSS 0.0476268f
c4 5 VSS 0.00503119f
c5 6 VSS 0.0041472f
c6 7 VSS 0.0046097f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1980 $X2=0.2970 $Y2=0.1665
r2 6 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1080 $X2=0.2970 $Y2=0.1215
r3 4 16 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r4 5 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r5 5 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1215
r6 5 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1665
r7 14 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r8 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r9 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r10 10 12 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r11 9 10 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r12 1 9 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r13 1 11 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r14 3 9 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r15 3 11 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r16 3 12 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_25 VSS 1
c1 1 VSS 0.0425523f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_27 VSS 1
c1 1 VSS 0.0425668f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_29 VSS 1
c1 1 VSS 0.0423487f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_28 VSS 1
c1 1 VSS 0.0423016f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_26 VSS 1
c1 1 VSS 0.0419712f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00521566f
.ends

.subckt PM_AND5x2_ASAP7_75t_R%NET14 VSS 21 22 83 86 88 90 92 94 96 3 29 24 4 5
+ 25 26 8 6 23 27 31 32 7 28 34 35 30 36 1 33
c1 1 VSS 0.0110556f
c2 3 VSS 0.00946489f
c3 4 VSS 0.00834735f
c4 5 VSS 0.00847044f
c5 6 VSS 0.00856271f
c6 7 VSS 0.00479636f
c7 8 VSS 0.00795894f
c8 21 VSS 0.0804992f
c9 22 VSS 0.08077f
c10 23 VSS 0.0024418f
c11 24 VSS 0.00464188f
c12 25 VSS 0.00475617f
c13 26 VSS 0.00411451f
c14 27 VSS 0.00429755f
c15 28 VSS 0.00385184f
c16 29 VSS 0.0731085f
c17 30 VSS 0.0133187f
c18 31 VSS 0.00346066f
c19 32 VSS 0.00385113f
c20 33 VSS 0.00125725f
c21 34 VSS 0.00315937f
c22 35 VSS 0.000450099f
c23 36 VSS 0.00362578f
r1 24 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r2 96 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r3 94 93 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r4 25 93 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r5 92 91 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 26 91 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 90 89 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r8 27 89 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.2025 $X2=0.6085 $Y2=0.2025
r9 88 87 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r10 28 87 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.2025 $X2=0.7705 $Y2=0.2025
r11 86 85 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7730 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r12 7 85 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7580 $Y=0.0675 $X2=0.7705 $Y2=0.0675
r13 82 7 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7460 $Y=0.0675 $X2=0.7580 $Y2=0.0675
r14 23 82 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7415 $Y=0.0675 $X2=0.7460 $Y2=0.0675
r15 83 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7390 $Y=0.0675 $X2=0.7415 $Y2=0.0675
r16 3 80 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.2340
r17 4 75 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2740 $Y2=0.2340
r18 5 73 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r19 6 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5980 $Y2=0.2340
r20 8 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.2025
+ $X2=0.7520 $Y2=0.2340
r21 7 58 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7560 $Y=0.0675
+ $X2=0.7560 $Y2=0.0360
r22 80 81 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.2135 $Y2=0.2340
r23 77 78 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2650 $Y2=0.2340
r24 77 81 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2135 $Y2=0.2340
r25 75 76 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.2340 $X2=0.2925 $Y2=0.2340
r26 75 78 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.2340 $X2=0.2650 $Y2=0.2340
r27 73 74 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r28 72 73 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r29 72 76 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.2925 $Y2=0.2340
r30 71 74 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4685
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r31 70 71 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4935
+ $Y=0.2340 $X2=0.4685 $Y2=0.2340
r32 69 70 10.8433 $w=1.3e-08 $l=4.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.4935 $Y2=0.2340
r33 67 68 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.2340 $X2=0.5890 $Y2=0.2340
r34 67 69 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r35 65 66 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5980
+ $Y=0.2340 $X2=0.6165 $Y2=0.2340
r36 65 68 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5980
+ $Y=0.2340 $X2=0.5890 $Y2=0.2340
r37 64 66 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.2340 $X2=0.6165 $Y2=0.2340
r38 62 63 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7335
+ $Y=0.2340 $X2=0.7520 $Y2=0.2340
r39 62 64 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7335
+ $Y=0.2340 $X2=0.6750 $Y2=0.2340
r40 60 61 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7610
+ $Y=0.2340 $X2=0.7945 $Y2=0.2340
r41 60 63 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.7610
+ $Y=0.2340 $X2=0.7520 $Y2=0.2340
r42 29 36 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8530 $Y=0.2340 $X2=0.8910 $Y2=0.2340
r43 29 61 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.8530
+ $Y=0.2340 $X2=0.7945 $Y2=0.2340
r44 58 59 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7560
+ $Y=0.0360 $X2=0.7945 $Y2=0.0360
r45 30 34 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8530 $Y=0.0360 $X2=0.8910 $Y2=0.0360
r46 30 59 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.8530
+ $Y=0.0360 $X2=0.7945 $Y2=0.0360
r47 36 56 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.2340 $X2=0.8910 $Y2=0.2160
r48 34 54 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0360 $X2=0.8910 $Y2=0.0540
r49 55 56 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1980 $X2=0.8910 $Y2=0.2160
r50 32 35 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.1665 $X2=0.8910 $Y2=0.1350
r51 32 55 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1665 $X2=0.8910 $Y2=0.1980
r52 53 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0720 $X2=0.8910 $Y2=0.0540
r53 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.0900 $X2=0.8910 $Y2=0.0720
r54 51 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1080 $X2=0.8910 $Y2=0.0900
r55 31 35 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.8910 $Y=0.1215 $X2=0.8910 $Y2=0.1350
r56 31 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.8910
+ $Y=0.1215 $X2=0.8910 $Y2=0.1080
r57 22 46 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.9990
+ $Y=0.1350 $X2=0.9990 $Y2=0.1350
r58 33 48 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.9095
+ $Y=0.1350 $X2=0.9280 $Y2=0.1350
r59 33 35 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.9095 $Y=0.1350 $X2=0.8910 $Y2=0.1350
r60 44 46 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9865 $Y=0.1350 $X2=0.9990 $Y2=0.1350
r61 43 44 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9720 $Y=0.1350 $X2=0.9865 $Y2=0.1350
r62 42 43 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.9575 $Y=0.1350 $X2=0.9720 $Y2=0.1350
r63 41 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.9245 $Y=0.1350
+ $X2=0.9280 $Y2=0.1350
r64 39 41 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.9325
+ $Y=0.1350 $X2=0.9245 $Y2=0.1350
r65 1 38 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.9360
+ $Y=0.1350 $X2=0.9460 $Y2=0.1350
r66 1 39 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.9360 $Y=0.1350 $X2=0.9325 $Y2=0.1350
r67 21 38 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9460 $Y2=0.1350
r68 21 39 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9325 $Y2=0.1350
r69 21 42 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.9450 $Y=0.1350 $X2=0.9575 $Y2=0.1350
r70 4 25 1e-05
r71 5 26 1e-05
r72 6 27 1e-05
r73 8 28 1e-05
.ends

.subckt PM_AND5x2_ASAP7_75t_R%C VSS 18 3 4 1 7 6
c1 1 VSS 0.00992208f
c2 3 VSS 0.00947513f
c3 4 VSS 0.0465653f
c4 5 VSS 0.00509654f
c5 6 VSS 0.00459911f
c6 7 VSS 0.00536955f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1980 $X2=0.4590 $Y2=0.1665
r2 3 15 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r3 18 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1665
r4 18 5 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1215
r5 5 6 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1215 $X2=0.4590 $Y2=0.1080
r6 13 15 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r7 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r8 11 12 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r9 10 17 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.4685
+ $Y=0.1350 $X2=0.4695 $Y2=0.1350
r10 9 10 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4685 $Y2=0.1350
r11 18 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1350
r12 1 9 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4495
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r13 1 11 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4495 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r14 4 9 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r15 4 11 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r16 4 17 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4695 $Y2=0.1350
.ends

.subckt PM_AND5x2_ASAP7_75t_R%NET35 VSS 11 14 22 25 1 7 2 8 9
c1 1 VSS 0.00478467f
c2 2 VSS 0.00491213f
c3 7 VSS 0.00228381f
c4 8 VSS 0.00226311f
c5 9 VSS 0.0213415f
r1 25 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r2 23 24 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6580 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r3 2 23 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6460 $Y=0.0675 $X2=0.6580 $Y2=0.0675
r4 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6460 $Y2=0.0675
r5 22 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
r6 2 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r7 18 19 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.6095
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r8 17 18 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.6095 $Y2=0.0360
r9 16 17 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4705
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r10 15 16 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4705 $Y2=0.0360
r11 9 15 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r12 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r13 14 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r14 1 13 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4340 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r15 10 1 0.148148 $w=8.1e-08 $l=1.2e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4220 $Y=0.0675 $X2=0.4340 $Y2=0.0675
r16 7 10 0.0555556 $w=8.1e-08 $l=4.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4220 $Y2=0.0675
r17 11 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
.ends

.subckt PM_AND5x2_ASAP7_75t_R%NET34 VSS 15 30 31 33 1 2 10 13 11 3 12
c1 1 VSS 0.00415771f
c2 2 VSS 0.00362746f
c3 3 VSS 0.00426633f
c4 10 VSS 0.00337691f
c5 11 VSS 0.00224181f
c6 12 VSS 0.00339158f
c7 13 VSS 0.00430739f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r3 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r4 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r6 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r7 3 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4820 $Y2=0.0720
r8 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0720
r9 24 25 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4635
+ $Y=0.0720 $X2=0.4820 $Y2=0.0720
r10 23 24 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4340
+ $Y=0.0720 $X2=0.4635 $Y2=0.0720
r11 22 23 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4025
+ $Y=0.0720 $X2=0.4340 $Y2=0.0720
r12 21 22 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0720 $X2=0.4025 $Y2=0.0720
r13 20 21 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3535
+ $Y=0.0720 $X2=0.3780 $Y2=0.0720
r14 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.0720 $X2=0.3535 $Y2=0.0720
r15 18 19 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2925
+ $Y=0.0720 $X2=0.3220 $Y2=0.0720
r16 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2740
+ $Y=0.0720 $X2=0.2925 $Y2=0.0720
r17 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2650
+ $Y=0.0720 $X2=0.2740 $Y2=0.0720
r18 13 16 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0720 $X2=0.2650 $Y2=0.0720
r19 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2740 $Y2=0.0720
r20 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r21 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r22 1 10 1e-05
.ends

.subckt PM_AND5x2_ASAP7_75t_R%NET32 VSS 15 30 31 33 1 2 10 13 11 3 12
c1 1 VSS 0.0038806f
c2 2 VSS 0.00321458f
c3 3 VSS 0.00417419f
c4 10 VSS 0.00301137f
c5 11 VSS 0.00207002f
c6 12 VSS 0.0029751f
c7 13 VSS 0.00365596f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7955 $Y=0.0675 $X2=0.8080 $Y2=0.0675
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7930 $Y=0.0675 $X2=0.7955 $Y2=0.0675
r3 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.7190 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r4 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.7020 $Y=0.0675 $X2=0.7165 $Y2=0.0675
r5 11 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6875 $Y=0.0675 $X2=0.7020 $Y2=0.0675
r6 30 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6850 $Y=0.0675 $X2=0.6875 $Y2=0.0675
r7 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.8100 $Y=0.0675
+ $X2=0.8100 $Y2=0.0720
r8 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.7020 $Y=0.0675
+ $X2=0.7020 $Y2=0.0720
r9 25 26 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.7790
+ $Y=0.0720 $X2=0.8100 $Y2=0.0720
r10 24 25 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.7495
+ $Y=0.0720 $X2=0.7790 $Y2=0.0720
r11 23 24 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.7310
+ $Y=0.0720 $X2=0.7495 $Y2=0.0720
r12 22 23 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.7155
+ $Y=0.0720 $X2=0.7310 $Y2=0.0720
r13 21 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.7020
+ $Y=0.0720 $X2=0.7155 $Y2=0.0720
r14 20 21 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.6775
+ $Y=0.0720 $X2=0.7020 $Y2=0.0720
r15 19 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6460
+ $Y=0.0720 $X2=0.6775 $Y2=0.0720
r16 18 19 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.6165
+ $Y=0.0720 $X2=0.6460 $Y2=0.0720
r17 17 18 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5980
+ $Y=0.0720 $X2=0.6165 $Y2=0.0720
r18 16 17 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5890
+ $Y=0.0720 $X2=0.5980 $Y2=0.0720
r19 13 16 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5825
+ $Y=0.0720 $X2=0.5890 $Y2=0.0720
r20 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5980 $Y2=0.0720
r21 15 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6110 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r22 10 14 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5960 $Y=0.0675 $X2=0.6085 $Y2=0.0675
r23 1 10 1e-05
.ends

.subckt PM_AND5x2_ASAP7_75t_R%B VSS 18 3 4 1 5 7 6
c1 1 VSS 0.012126f
c2 3 VSS 0.0461325f
c3 4 VSS 0.0476139f
c4 5 VSS 0.00509407f
c5 6 VSS 0.00447098f
c6 7 VSS 0.00487886f
r1 7 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1980 $X2=0.6210 $Y2=0.1665
r2 4 16 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r3 18 19 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1665
r4 18 5 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1215
r5 5 6 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1215 $X2=0.6210 $Y2=0.1080
r6 14 16 5.66664 $w=1.866e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6625 $Y=0.1350 $X2=0.6750 $Y2=0.1350
r7 13 14 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6480 $Y=0.1350 $X2=0.6625 $Y2=0.1350
r8 12 13 14.4473 $w=1.33e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.6335 $Y=0.1350 $X2=0.6480 $Y2=0.1350
r9 10 12 2.64971 $w=1.44167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.6305 $Y=0.1350 $X2=0.6335 $Y2=0.1350
r10 9 10 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6305 $Y2=0.1350
r11 18 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
r12 1 9 3.01694 $w=2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.6115
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r13 1 11 0.65697 $w=1.665e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.6115
+ $Y=0.1350 $X2=0.6105 $Y2=0.1350
r14 3 9 3.17282 $w=1.28947e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r15 3 11 0.812849 $w=2.16824e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6105 $Y2=0.1350
r16 3 12 2.80558 $w=1.8426e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.6210 $Y=0.1350 $X2=0.6335 $Y2=0.1350
.ends


*
.SUBCKT AND5x2_ASAP7_75t_R VSS VDD E D C B A Y
*
* VSS VSS
* VDD VDD
* E E
* D D
* C C
* B B
* A A
* Y Y
*
*

MM6 N_MM6_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM5@2_g N_MM5@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 N_MM3@2_d N_MM8_g N_MM3@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM7_g N_MM4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM10_g N_MM0@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM11@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "AND5x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "AND5x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_AND5x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_AND5x2_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM6_g 0.00247251f
x_PM_AND5x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_AND5x2_ASAP7_75t_R%noxref_15
cc_2 N_noxref_15_1 N_MM6_g 0.0104075f
cc_3 N_noxref_15_1 N_noxref_14_1 0.00193994f
x_PM_AND5x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_AND5x2_ASAP7_75t_R%noxref_18
cc_4 N_noxref_18_1 N_MM2_g 0.00146234f
cc_5 N_noxref_18_1 N_NET34_10 0.0357044f
cc_6 N_noxref_18_1 N_noxref_16_1 0.00766796f
x_PM_AND5x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_AND5x2_ASAP7_75t_R%noxref_16
cc_7 N_noxref_16_1 N_MM9_g 0.0013953f
cc_8 N_noxref_16_1 N_NET34_10 0.000580909f
x_PM_AND5x2_ASAP7_75t_R%NET33 VSS N_MM6_d N_MM6@2_d N_MM5_s N_MM5@2_s N_NET33_1
+ N_NET33_7 N_NET33_2 N_NET33_8 N_NET33_9 PM_AND5x2_ASAP7_75t_R%NET33
cc_9 N_NET33_1 N_MM6_g 0.00196267f
cc_10 N_NET33_7 N_E_1 0.00209113f
cc_11 N_NET33_7 N_MM9_g 0.0182001f
cc_12 N_NET33_7 N_MM6_g 0.0505108f
cc_13 N_NET33_2 N_MM2_g 0.00188663f
cc_14 N_NET33_8 N_D_1 0.0019024f
cc_15 N_NET33_8 N_MM5@2_g 0.0182102f
cc_16 N_NET33_8 N_MM2_g 0.049378f
x_PM_AND5x2_ASAP7_75t_R%noxref_22 VSS N_noxref_22_1
+ PM_AND5x2_ASAP7_75t_R%noxref_22
cc_17 N_noxref_22_1 N_MM7_g 0.00144396f
cc_18 N_noxref_22_1 N_NET34_12 0.000574837f
cc_19 N_noxref_22_1 N_NET32_10 0.0355455f
cc_20 N_noxref_22_1 N_noxref_20_1 0.00766795f
x_PM_AND5x2_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1
+ PM_AND5x2_ASAP7_75t_R%noxref_20
cc_21 N_noxref_20_1 N_MM8_g 0.0014579f
cc_22 N_noxref_20_1 N_NET34_12 0.0359828f
cc_23 N_noxref_20_1 N_NET32_10 0.000574573f
x_PM_AND5x2_ASAP7_75t_R%noxref_23 VSS N_noxref_23_1
+ PM_AND5x2_ASAP7_75t_R%noxref_23
cc_24 N_noxref_23_1 N_MM7_g 0.00148184f
cc_25 N_noxref_23_1 N_NET14_6 0.000422069f
cc_26 N_noxref_23_1 N_NET14_27 0.0368478f
cc_27 N_noxref_23_1 N_noxref_21_1 0.00765415f
cc_28 N_noxref_23_1 N_noxref_22_1 0.00123971f
x_PM_AND5x2_ASAP7_75t_R%Y VSS Y N_MM11_d N_MM11@2_d N_MM1_d N_MM1@2_d N_Y_7
+ N_Y_2 N_Y_8 N_Y_11 N_Y_1 PM_AND5x2_ASAP7_75t_R%Y
cc_29 N_Y_7 N_NET14_29 0.000101606f
cc_30 N_Y_7 N_NET14_34 0.000161247f
cc_31 N_Y_7 N_NET14_36 0.000174871f
cc_32 N_Y_7 N_NET14_1 0.000425186f
cc_33 N_Y_7 N_NET14_31 0.000499674f
cc_34 N_Y_7 N_NET14_32 0.000511823f
cc_35 N_Y_7 N_MM11@2_g 0.0384511f
cc_36 N_Y_2 N_NET14_33 0.000664079f
cc_37 N_Y_8 N_MM11_g 0.0311268f
cc_38 N_Y_11 N_NET14_1 0.000890406f
cc_39 N_Y_1 N_MM11_g 0.00204472f
cc_40 N_Y_2 N_MM11_g 0.00214898f
cc_41 N_Y_8 N_NET14_1 0.00490255f
cc_42 N_Y_7 N_MM11_g 0.0690454f
x_PM_AND5x2_ASAP7_75t_R%A VSS A N_MM0_g N_MM10_g N_A_5 N_A_1 N_A_7 N_A_6
+ PM_AND5x2_ASAP7_75t_R%A
cc_43 N_MM0_g N_B_1 0.00141624f
cc_44 N_MM0_g N_MM4@2_g 0.0124892f
x_PM_AND5x2_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1
+ PM_AND5x2_ASAP7_75t_R%noxref_21
cc_45 N_noxref_21_1 N_MM8_g 0.00149404f
cc_46 N_noxref_21_1 N_NET14_6 0.000138562f
cc_47 N_noxref_21_1 N_NET14_26 0.000632803f
cc_48 N_noxref_21_1 N_noxref_20_1 0.00124092f
x_PM_AND5x2_ASAP7_75t_R%E VSS E N_MM6_g N_MM9_g N_E_1 PM_AND5x2_ASAP7_75t_R%E
x_PM_AND5x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_AND5x2_ASAP7_75t_R%noxref_17
cc_49 N_noxref_17_1 N_MM9_g 0.00139123f
cc_50 N_noxref_17_1 N_NET14_4 0.000140192f
cc_51 N_noxref_17_1 N_NET14_3 0.00043218f
cc_52 N_noxref_17_1 N_NET14_24 0.0369805f
cc_53 N_noxref_17_1 N_noxref_16_1 0.00123565f
x_PM_AND5x2_ASAP7_75t_R%noxref_24 VSS N_noxref_24_1
+ PM_AND5x2_ASAP7_75t_R%noxref_24
cc_54 N_noxref_24_1 N_MM10_g 0.00139398f
cc_55 N_noxref_24_1 N_NET14_23 0.000537822f
cc_56 N_noxref_24_1 N_NET32_12 0.0358517f
x_PM_AND5x2_ASAP7_75t_R%D VSS D N_MM2_g N_MM5@2_g N_D_1 N_D_7 N_D_6
+ PM_AND5x2_ASAP7_75t_R%D
x_PM_AND5x2_ASAP7_75t_R%noxref_25 VSS N_noxref_25_1
+ PM_AND5x2_ASAP7_75t_R%noxref_25
cc_57 N_noxref_25_1 N_MM10_g 0.00141569f
cc_58 N_noxref_25_1 N_NET14_32 7.26266e-20
cc_59 N_noxref_25_1 N_NET14_28 0.00047975f
cc_60 N_noxref_25_1 N_noxref_24_1 0.00123888f
x_PM_AND5x2_ASAP7_75t_R%noxref_27 VSS N_noxref_27_1
+ PM_AND5x2_ASAP7_75t_R%noxref_27
cc_61 N_noxref_27_1 N_NET14_32 8.51408e-20
cc_62 N_noxref_27_1 N_MM11_g 0.00179085f
cc_63 N_noxref_27_1 N_noxref_25_1 0.00764661f
cc_64 N_noxref_27_1 N_noxref_26_1 0.00121702f
x_PM_AND5x2_ASAP7_75t_R%noxref_29 VSS N_noxref_29_1
+ PM_AND5x2_ASAP7_75t_R%noxref_29
cc_65 N_noxref_29_1 N_MM11@2_g 0.00145483f
cc_66 N_noxref_29_1 N_Y_8 0.000854864f
cc_67 N_noxref_29_1 N_noxref_28_1 0.00176693f
x_PM_AND5x2_ASAP7_75t_R%noxref_28 VSS N_noxref_28_1
+ PM_AND5x2_ASAP7_75t_R%noxref_28
cc_68 N_noxref_28_1 N_MM11@2_g 0.00145781f
cc_69 N_noxref_28_1 N_Y_7 0.000853981f
x_PM_AND5x2_ASAP7_75t_R%noxref_26 VSS N_noxref_26_1
+ PM_AND5x2_ASAP7_75t_R%noxref_26
cc_70 N_noxref_26_1 N_NET14_31 8.36024e-20
cc_71 N_noxref_26_1 N_MM11_g 0.00178625f
cc_72 N_noxref_26_1 N_NET32_12 0.000576438f
cc_73 N_noxref_26_1 N_noxref_24_1 0.00766318f
x_PM_AND5x2_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1
+ PM_AND5x2_ASAP7_75t_R%noxref_19
cc_74 N_noxref_19_1 N_MM2_g 0.0014903f
cc_75 N_noxref_19_1 N_NET14_3 0.000147408f
cc_76 N_noxref_19_1 N_NET14_4 0.000421868f
cc_77 N_noxref_19_1 N_NET14_25 0.0372598f
cc_78 N_noxref_19_1 N_noxref_17_1 0.00767868f
cc_79 N_noxref_19_1 N_noxref_18_1 0.00123876f
x_PM_AND5x2_ASAP7_75t_R%NET14 VSS N_MM11_g N_MM11@2_g N_MM0_d N_MM0@2_d
+ N_MM10_d N_MM7_d N_MM8_d N_MM2_d N_MM9_d N_NET14_3 N_NET14_29 N_NET14_24
+ N_NET14_4 N_NET14_5 N_NET14_25 N_NET14_26 N_NET14_8 N_NET14_6 N_NET14_23
+ N_NET14_27 N_NET14_31 N_NET14_32 N_NET14_7 N_NET14_28 N_NET14_34 N_NET14_35
+ N_NET14_30 N_NET14_36 N_NET14_1 N_NET14_33 PM_AND5x2_ASAP7_75t_R%NET14
cc_80 N_NET14_3 N_MM9_g 0.00131589f
cc_81 N_NET14_29 N_MM9_g 0.000536096f
cc_82 N_NET14_24 N_E_1 0.00102901f
cc_83 N_NET14_24 N_MM9_g 0.0349314f
cc_84 N_NET14_3 N_MM2_g 0.000114593f
cc_85 N_NET14_4 N_MM2_g 0.0026646f
cc_86 N_NET14_5 N_MM2_g 0.000237021f
cc_87 N_NET14_4 N_D 0.000957312f
cc_88 N_NET14_25 N_D_1 0.00101646f
cc_89 N_NET14_29 N_D_7 0.00589377f
cc_90 N_NET14_25 N_MM2_g 0.0357843f
cc_91 N_NET14_5 N_MM3_g 0.00413968f
cc_92 N_NET14_26 N_MM8_g 0.0310845f
cc_93 N_NET14_26 N_C_1 0.00235505f
cc_94 N_NET14_29 N_MM3_g 0.00263317f
cc_95 N_NET14_29 N_C_7 0.00291898f
cc_96 N_NET14_26 N_MM3_g 0.0411297f
cc_97 N_NET14_8 N_MM7_g 0.00016563f
cc_98 N_NET14_6 N_MM7_g 0.00253496f
cc_99 N_NET14_23 N_MM7_g 0.000380076f
cc_100 N_NET14_6 N_B_5 0.000952829f
cc_101 N_NET14_27 N_B_1 0.00103653f
cc_102 N_NET14_29 N_B_7 0.00540195f
cc_103 N_NET14_27 N_MM7_g 0.0354082f
cc_104 N_NET14_31 N_MM0_g 0.000132739f
cc_105 N_NET14_32 N_MM0_g 0.000170113f
cc_106 N_NET14_8 N_MM0_g 0.00355667f
cc_107 N_NET14_7 N_MM0_g 0.00256455f
cc_108 N_NET14_8 N_A_5 0.00110754f
cc_109 N_NET14_28 N_MM10_g 0.0123281f
cc_110 N_NET14_28 N_A_1 0.00435607f
cc_111 N_NET14_29 N_A_7 0.00585776f
cc_112 N_NET14_28 N_MM0_g 0.0214932f
cc_113 N_NET14_23 N_MM10_g 0.0379342f
cc_114 N_NET14_23 N_MM0_g 0.0701759f
x_PM_AND5x2_ASAP7_75t_R%C VSS C N_MM3_g N_MM8_g N_C_1 N_C_7 N_C_6
+ PM_AND5x2_ASAP7_75t_R%C
cc_115 N_MM3_g N_MM5@2_g 0.0128576f
x_PM_AND5x2_ASAP7_75t_R%NET35 VSS N_MM3_d N_MM3@2_d N_MM4_s N_MM4@2_s N_NET35_1
+ N_NET35_7 N_NET35_2 N_NET35_8 N_NET35_9 PM_AND5x2_ASAP7_75t_R%NET35
cc_116 N_NET35_1 N_MM3_g 0.00188569f
cc_117 N_NET35_7 N_C_1 0.00190001f
cc_118 N_NET35_7 N_MM8_g 0.0181683f
cc_119 N_NET35_7 N_MM3_g 0.049176f
cc_120 N_NET35_2 N_MM7_g 0.00188077f
cc_121 N_NET35_8 N_B_1 0.00202515f
cc_122 N_NET35_8 N_MM4@2_g 0.0181993f
cc_123 N_NET35_8 N_MM7_g 0.0492077f
cc_124 N_NET35_9 N_NET34_12 0.000594811f
cc_125 N_NET35_1 N_NET34_13 0.000744847f
cc_126 N_NET35_7 N_NET34_11 0.00112085f
cc_127 N_NET35_1 N_NET34_3 0.00173686f
cc_128 N_NET35_1 N_NET34_2 0.00434073f
cc_129 N_NET35_9 N_NET34_13 0.0101514f
x_PM_AND5x2_ASAP7_75t_R%NET34 VSS N_MM5_d N_MM5@2_d N_MM3_s N_MM3@2_s N_NET34_1
+ N_NET34_2 N_NET34_10 N_NET34_13 N_NET34_11 N_NET34_3 N_NET34_12
+ PM_AND5x2_ASAP7_75t_R%NET34
cc_130 N_NET34_1 N_MM5@2_g 0.000576559f
cc_131 N_NET34_2 N_MM5@2_g 0.000759812f
cc_132 N_NET34_1 N_MM2_g 0.00116896f
cc_133 N_NET34_10 N_D_1 0.0017025f
cc_134 N_NET34_13 N_D_6 0.00521131f
cc_135 N_NET34_10 N_MM2_g 0.0333262f
cc_136 N_NET34_11 N_MM5@2_g 0.0350704f
cc_137 N_NET34_2 N_MM3_g 0.000777644f
cc_138 N_NET34_3 N_MM8_g 0.00114437f
cc_139 N_NET34_11 N_C_1 0.00170317f
cc_140 N_NET34_13 N_C_6 0.00512374f
cc_141 N_NET34_11 N_MM3_g 0.0332558f
cc_142 N_NET34_12 N_MM8_g 0.0356687f
cc_143 N_NET34_10 N_NET33_9 0.000604248f
cc_144 N_NET34_10 N_NET33_8 0.00112311f
cc_145 N_NET34_2 N_NET33_2 0.0012574f
cc_146 N_NET34_1 N_NET33_2 0.00485848f
cc_147 N_NET34_13 N_NET33_9 0.0110467f
x_PM_AND5x2_ASAP7_75t_R%NET32 VSS N_MM4_d N_MM4@2_d N_MM0_s N_MM0@2_s N_NET32_1
+ N_NET32_2 N_NET32_10 N_NET32_13 N_NET32_11 N_NET32_3 N_NET32_12
+ PM_AND5x2_ASAP7_75t_R%NET32
cc_148 N_NET32_1 N_MM4@2_g 0.000477502f
cc_149 N_NET32_2 N_MM4@2_g 0.000745474f
cc_150 N_NET32_1 N_MM7_g 0.00114406f
cc_151 N_NET32_10 N_B_1 0.00173373f
cc_152 N_NET32_13 N_B_6 0.0047129f
cc_153 N_NET32_10 N_MM7_g 0.0331856f
cc_154 N_NET32_11 N_MM4@2_g 0.0349308f
cc_155 N_NET32_2 N_MM0_g 0.0015514f
cc_156 N_NET32_3 N_MM0_g 0.000858279f
cc_157 N_NET32_11 N_A_1 0.00167693f
cc_158 N_NET32_13 N_A_6 0.00490804f
cc_159 N_NET32_12 N_MM10_g 0.0331987f
cc_160 N_NET32_11 N_MM0_g 0.0349173f
cc_161 N_NET32_13 N_NET14_8 4.67999e-20
cc_162 N_NET32_13 N_NET14_27 0.000415716f
cc_163 N_NET32_13 N_NET14_34 5.73913e-20
cc_164 N_NET32_13 N_NET14_23 0.000101698f
cc_165 N_NET32_13 N_NET14_32 0.00015872f
cc_166 N_NET32_13 N_NET14_6 0.000160867f
cc_167 N_NET32_13 N_NET14_35 0.000161268f
cc_168 N_NET32_13 N_NET14_29 0.000226391f
cc_169 N_NET32_2 N_NET14_7 0.00456101f
cc_170 N_NET32_13 N_NET14_31 0.000550033f
cc_171 N_NET32_11 N_NET14_23 0.00169266f
cc_172 N_NET32_12 N_NET14_23 0.000652875f
cc_173 N_NET32_13 N_NET14_7 0.000694971f
cc_174 N_NET32_3 N_NET14_30 0.00089415f
cc_175 N_NET32_3 N_NET14_7 0.00202246f
cc_176 N_NET32_13 N_NET14_30 0.0094372f
cc_177 N_NET32_1 N_NET35_9 0.000597982f
cc_178 N_NET32_13 N_NET35_2 0.000822453f
cc_179 N_NET32_10 N_NET35_8 0.00112157f
cc_180 N_NET32_2 N_NET35_2 0.00126176f
cc_181 N_NET32_1 N_NET35_2 0.00479583f
cc_182 N_NET32_13 N_NET35_9 0.0101298f
x_PM_AND5x2_ASAP7_75t_R%B VSS B N_MM7_g N_MM4@2_g N_B_1 N_B_5 N_B_7 N_B_6
+ PM_AND5x2_ASAP7_75t_R%B
*END of AND5x2_ASAP7_75t_R.pxi
.ENDS
** Design:	OR2x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR2x2_ASAP7_75t_R%NET15 VSS 2 3 1
c1 1 VSS 0.000951754f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR2x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0423665f
.ends

.subckt PM_OR2x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0423633f
.ends

.subckt PM_OR2x2_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0048651f
.ends

.subckt PM_OR2x2_ASAP7_75t_R%B VSS 18 3 1 6 7 5
c1 1 VSS 0.00186336f
c2 3 VSS 0.0328897f
c3 4 VSS 0.0071564f
c4 5 VSS 0.0051706f
c5 6 VSS 0.00167966f
c6 7 VSS 0.00783327f
c7 8 VSS 0.00159643f
r1 7 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 5 19 5.73148 $w=1.38716e-08 $l=2.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1392
r3 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r4 4 8 5.62944 $w=1.37143e-08 $l=2.62e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1297
r5 4 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r6 18 19 0.535733 $w=1.8e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1340 $X2=0.0270 $Y2=0.1392
r7 18 8 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1340 $X2=0.0270 $Y2=0.1297
r8 18 15 0.517402 $w=3.18182e-09 $l=1.10454e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1340 $X2=0.0380 $Y2=0.1350
r9 14 16 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0545
+ $Y=0.1350 $X2=0.0635 $Y2=0.1350
r10 6 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0470
+ $Y=0.1350 $X2=0.0545 $Y2=0.1350
r11 6 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0470
+ $Y=0.1350 $X2=0.0380 $Y2=0.1350
r12 12 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0600 $Y=0.1355
+ $X2=0.0635 $Y2=0.1350
r13 11 12 3.89665 $w=1.63e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0685 $Y=0.1355 $X2=0.0600 $Y2=0.1355
r14 1 10 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1355 $X2=0.0815 $Y2=0.1355
r15 1 11 1.26439 $w=1.74167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0715 $Y=0.1355 $X2=0.0685 $Y2=0.1355
r16 3 10 2.56268 $w=1.27615e-07 $l=7.07107e-10 $layer=LIG
+ $thickness=5.21026e-08 $X=0.0810 $Y=0.1350 $X2=0.0815 $Y2=0.1355
r17 3 11 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1355
.ends

.subckt PM_OR2x2_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0315713f
.ends

.subckt PM_OR2x2_ASAP7_75t_R%Y VSS 28 20 21 36 37 7 1 13 9 14 15 2 10 8
c1 1 VSS 0.00861159f
c2 2 VSS 0.00856141f
c3 7 VSS 0.00463849f
c4 8 VSS 0.00456362f
c5 9 VSS 0.00125944f
c6 10 VSS 0.00102072f
c7 11 VSS 0.00656615f
c8 12 VSS 0.00666974f
c9 13 VSS 0.00741181f
c10 14 VSS 0.00225515f
c11 15 VSS 0.00273782f
c12 16 VSS 0.00351869f
c13 17 VSS 0.00350735f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 36 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2160 $Y2=0.2160
r7 10 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1865 $X2=0.2160 $Y2=0.1980
r8 15 31 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2260 $Y2=0.2340
r9 15 33 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2160 $Y2=0.2160
r10 12 17 7.56188 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2575 $Y=0.2340 $X2=0.2970 $Y2=0.2340
r11 12 31 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2575
+ $Y=0.2340 $X2=0.2260 $Y2=0.2340
r12 17 30 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.2340 $X2=0.2970 $Y2=0.2045
r13 29 30 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1660 $X2=0.2970 $Y2=0.2045
r14 28 29 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1660
r15 28 27 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1455
r16 26 27 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1455
r17 25 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1060 $X2=0.2970 $Y2=0.1350
r18 13 16 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0655 $X2=0.2970 $Y2=0.0360
r19 13 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0655 $X2=0.2970 $Y2=0.1060
r20 16 24 7.56188 $w=1.41392e-08 $l=3.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2575 $Y2=0.0360
r21 11 14 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2260
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r22 11 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2260
+ $Y=0.0360 $X2=0.2575 $Y2=0.0360
r23 9 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0720
r24 9 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0360
r25 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r26 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r27 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r28 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r29 20 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends

.subckt PM_OR2x2_ASAP7_75t_R%A VSS 4 3 1 5 6
c1 1 VSS 0.00553121f
c2 3 VSS 0.082582f
c3 4 VSS 0.00263751f
c4 5 VSS 0.00188427f
c5 6 VSS 0.00189829f
r1 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 9 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r4 4 10 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1665
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_OR2x2_ASAP7_75t_R%NET7 VSS 9 10 53 54 56 14 3 4 13 12 11 19 1 15 16
+ 17 18 20
c1 1 VSS 0.0070048f
c2 3 VSS 0.007042f
c3 4 VSS 0.00923767f
c4 9 VSS 0.0805255f
c5 10 VSS 0.0807903f
c6 11 VSS 0.00691717f
c7 12 VSS 0.00659148f
c8 13 VSS 0.0143804f
c9 14 VSS 0.00867471f
c10 15 VSS 0.00274963f
c11 16 VSS 0.00272149f
c12 17 VSS 0.0011368f
c13 18 VSS 0.00221803f
c14 19 VSS 0.000164379f
c15 20 VSS 0.00257171f
r1 56 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 12 55 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 54 52 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r4 4 52 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r5 11 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r6 53 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r7 3 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r8 4 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1120 $Y2=0.0360
r9 49 50 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0700 $Y2=0.2340
r10 47 50 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.2340 $X2=0.0700 $Y2=0.2340
r11 46 47 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1005
+ $Y=0.2340 $X2=0.0855 $Y2=0.2340
r12 45 46 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1005 $Y2=0.2340
r13 13 20 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1560 $Y=0.2340 $X2=0.1770 $Y2=0.2340
r14 13 45 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1560
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r15 41 42 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r16 14 18 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1560 $Y=0.0360 $X2=0.1770 $Y2=0.0360
r17 14 42 5.94634 $w=1.3e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1560
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r18 20 40 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.2340 $X2=0.1770 $Y2=0.2160
r19 18 37 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.0360 $X2=0.1770 $Y2=0.0540
r20 39 40 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.1980 $X2=0.1770 $Y2=0.2160
r21 38 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.1865 $X2=0.1770 $Y2=0.1980
r22 16 19 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1770 $Y=0.1640 $X2=0.1770 $Y2=0.1350
r23 16 38 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.1640 $X2=0.1770 $Y2=0.1865
r24 36 37 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.0720 $X2=0.1770 $Y2=0.0540
r25 35 36 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.0835 $X2=0.1770 $Y2=0.0720
r26 15 19 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1770 $Y=0.1060 $X2=0.1770 $Y2=0.1350
r27 15 35 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.1060 $X2=0.1770 $Y2=0.0835
r28 10 28 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r29 30 31 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2055
+ $Y=0.1350 $X2=0.2145 $Y2=0.1350
r30 17 30 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1950
+ $Y=0.1350 $X2=0.2055 $Y2=0.1350
r31 17 19 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1950
+ $Y=0.1350 $X2=0.1770 $Y2=0.1350
r32 26 28 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r33 25 26 3.24898 $w=1.53e-08 $l=5.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2250 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r34 24 25 7.08868 $w=1.53e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2130 $Y=0.1350 $X2=0.2250 $Y2=0.1350
r35 24 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2130 $Y=0.1350
+ $X2=0.2145 $Y2=0.1350
r36 23 24 6.79332 $w=1.53e-08 $l=1.15e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.2130 $Y2=0.1350
r37 9 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r38 1 22 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r39 1 23 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r40 9 22 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r41 9 23 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r42 3 12 1e-05
.ends


*
.SUBCKT OR2x2_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 VSS N_MM5_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 VSS N_MM5@2_g N_MM5@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM2_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VDD N_MM5_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 VDD N_MM5@2_g N_MM0@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR2x2_ASAP7_75t_R%NET15 VSS N_MM4_d N_MM3_s N_NET15_1
+ PM_OR2x2_ASAP7_75t_R%NET15
cc_1 N_NET15_1 N_MM1_g 0.0173983f
cc_2 N_NET15_1 N_MM2_g 0.0173768f
x_PM_OR2x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR2x2_ASAP7_75t_R%noxref_11
cc_3 N_noxref_11_1 N_MM5@2_g 0.00147549f
cc_4 N_noxref_11_1 N_Y_8 0.000845022f
cc_5 N_noxref_11_1 N_noxref_10_1 0.00177919f
x_PM_OR2x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR2x2_ASAP7_75t_R%noxref_10
cc_6 N_noxref_10_1 N_MM5@2_g 0.00146996f
cc_7 N_noxref_10_1 N_Y_7 0.000846712f
x_PM_OR2x2_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_OR2x2_ASAP7_75t_R%noxref_9
cc_8 N_noxref_9_1 N_MM1_g 0.00249476f
cc_9 N_noxref_9_1 N_NET7_12 0.0372529f
cc_10 N_noxref_9_1 N_noxref_8_1 0.00186f
x_PM_OR2x2_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_6 N_B_7 N_B_5
+ PM_OR2x2_ASAP7_75t_R%B
x_PM_OR2x2_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1 PM_OR2x2_ASAP7_75t_R%noxref_8
cc_11 N_noxref_8_1 N_MM1_g 0.00467413f
cc_12 N_noxref_8_1 N_NET7_11 0.000579783f
x_PM_OR2x2_ASAP7_75t_R%Y VSS Y N_MM5_s N_MM5@2_s N_MM0_s N_MM0@2_s N_Y_7 N_Y_1
+ N_Y_13 N_Y_9 N_Y_14 N_Y_15 N_Y_2 N_Y_10 N_Y_8 PM_OR2x2_ASAP7_75t_R%Y
cc_13 N_Y_7 N_NET7_16 0.00060676f
cc_14 N_Y_1 N_NET7_1 0.000989123f
cc_15 N_Y_13 N_NET7_1 0.00103517f
cc_16 N_Y_9 N_NET7_17 0.0013171f
cc_17 N_Y_14 N_NET7_18 0.00146395f
cc_18 N_Y_15 N_NET7_20 0.00146468f
cc_19 N_Y_1 N_MM5@2_g 0.0022066f
cc_20 N_Y_2 N_MM5@2_g 0.00220838f
cc_21 N_Y_9 N_NET7_15 0.00402762f
cc_22 N_Y_10 N_NET7_16 0.00405057f
cc_23 N_Y_8 N_NET7_1 0.00455125f
cc_24 N_Y_8 N_MM5@2_g 0.0302457f
cc_25 N_Y_7 N_MM5_g 0.0373798f
cc_26 N_Y_7 N_MM5@2_g 0.0707074f
x_PM_OR2x2_ASAP7_75t_R%A VSS A N_MM2_g N_A_1 N_A_5 N_A_6 PM_OR2x2_ASAP7_75t_R%A
cc_27 N_MM2_g N_B_1 0.000402027f
cc_28 N_MM2_g N_B_6 0.000490086f
cc_29 N_A_1 N_B_1 0.00175859f
cc_30 N_A N_B_6 0.00176934f
cc_31 N_MM2_g N_MM1_g 0.00841607f
x_PM_OR2x2_ASAP7_75t_R%NET7 VSS N_MM5_g N_MM5@2_g N_MM1_s N_MM2_s N_MM4_s
+ N_NET7_14 N_NET7_3 N_NET7_4 N_NET7_13 N_NET7_12 N_NET7_11 N_NET7_19 N_NET7_1
+ N_NET7_15 N_NET7_16 N_NET7_17 N_NET7_18 N_NET7_20 PM_OR2x2_ASAP7_75t_R%NET7
cc_32 N_NET7_14 N_MM1_g 0.000381532f
cc_33 N_NET7_3 N_B_6 0.000422175f
cc_34 N_NET7_3 N_B_1 0.000533292f
cc_35 N_NET7_4 N_MM1_g 0.000614776f
cc_36 N_NET7_14 N_B_7 0.000846721f
cc_37 N_NET7_13 N_B_5 0.000947128f
cc_38 N_NET7_3 N_B_5 0.00156148f
cc_39 N_NET7_12 N_B_1 0.00189624f
cc_40 N_NET7_3 N_MM1_g 0.00250821f
cc_41 N_NET7_11 N_MM1_g 0.0109883f
cc_42 N_NET7_12 N_MM1_g 0.0505924f
cc_43 N_NET7_3 N_MM2_g 0.000410267f
cc_44 N_NET7_19 N_MM2_g 0.000579268f
cc_45 N_NET7_4 N_MM2_g 0.000810524f
cc_46 N_NET7_1 N_A_1 0.00128577f
cc_47 N_NET7_15 N_A 0.00185829f
cc_48 N_NET7_16 N_A 0.00202616f
cc_49 N_NET7_11 N_MM2_g 0.0110302f
cc_50 N_NET7_19 N_A 0.00438262f
cc_51 N_NET7_14 N_A_5 0.00481714f
cc_52 N_NET7_13 N_A_6 0.00493847f
cc_53 N_MM5_g N_MM2_g 0.018311f
*END of OR2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	OR2x4_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR2x4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR2x4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR2x4_ASAP7_75t_R%NET15 VSS 2 3 1
c1 1 VSS 0.000951677f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR2x4_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0048411f
.ends

.subckt PM_OR2x4_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0315345f
.ends

.subckt PM_OR2x4_ASAP7_75t_R%A VSS 4 3 1 5 6
c1 1 VSS 0.00565419f
c2 3 VSS 0.0825559f
c3 4 VSS 0.00274027f
c4 5 VSS 0.00192312f
c5 6 VSS 0.00199917f
r1 6 10 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 5 9 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 9 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1035
r4 4 10 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1665
r5 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r6 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_OR2x4_ASAP7_75t_R%B VSS 18 3 6 1 7 5
c1 1 VSS 0.00194742f
c2 3 VSS 0.0329006f
c3 4 VSS 0.0071658f
c4 5 VSS 0.00515311f
c5 6 VSS 0.00167855f
c6 7 VSS 0.00786434f
c7 8 VSS 0.00161097f
r1 7 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r2 5 19 5.73148 $w=1.38716e-08 $l=2.73e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1392
r3 20 21 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r4 4 8 5.62944 $w=1.37143e-08 $l=2.62e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1297
r5 4 20 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r6 18 19 0.535733 $w=1.8e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1340 $X2=0.0270 $Y2=0.1392
r7 18 8 0.433689 $w=1.8e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1340 $X2=0.0270 $Y2=0.1297
r8 18 15 0.517402 $w=3.18182e-09 $l=1.10454e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1340 $X2=0.0380 $Y2=0.1350
r9 14 16 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0545
+ $Y=0.1350 $X2=0.0635 $Y2=0.1350
r10 6 14 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0470
+ $Y=0.1350 $X2=0.0545 $Y2=0.1350
r11 6 15 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0470
+ $Y=0.1350 $X2=0.0380 $Y2=0.1350
r12 12 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0600 $Y=0.1355
+ $X2=0.0635 $Y2=0.1350
r13 11 12 3.89665 $w=1.63e-08 $l=8.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0685 $Y=0.1355 $X2=0.0600 $Y2=0.1355
r14 1 10 2.36633 $w=2.3e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1355 $X2=0.0815 $Y2=0.1355
r15 1 11 1.26439 $w=1.74167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0715 $Y=0.1355 $X2=0.0685 $Y2=0.1355
r16 3 10 2.56268 $w=1.27615e-07 $l=7.07107e-10 $layer=LIG
+ $thickness=5.21026e-08 $X=0.0810 $Y=0.1350 $X2=0.0815 $Y2=0.1355
r17 3 11 1.46074 $w=1.8486e-07 $l=1.251e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1355
.ends

.subckt PM_OR2x4_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0422849f
.ends

.subckt PM_OR2x4_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0422849f
.ends

.subckt PM_OR2x4_ASAP7_75t_R%NET7 VSS 9 10 11 12 68 69 71 13 16 3 4 15 14 1 21
+ 17 18 22 20 19
c1 1 VSS 0.0188773f
c2 3 VSS 0.0086887f
c3 4 VSS 0.0116595f
c4 9 VSS 0.0816395f
c5 10 VSS 0.0815519f
c6 11 VSS 0.0813273f
c7 12 VSS 0.081932f
c8 13 VSS 0.00784891f
c9 14 VSS 0.00653321f
c10 15 VSS 0.0141053f
c11 16 VSS 0.00857084f
c12 17 VSS 0.003176f
c13 18 VSS 0.00322497f
c14 19 VSS 0.00202273f
c15 20 VSS 0.00401353f
c16 21 VSS 0.00142359f
c17 22 VSS 0.00383463f
r1 71 70 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 14 70 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 69 67 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r4 4 67 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r5 13 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r6 68 13 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r7 3 64 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r8 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1120 $Y2=0.0360
r9 64 65 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0700 $Y2=0.2340
r10 62 65 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0855
+ $Y=0.2340 $X2=0.0700 $Y2=0.2340
r11 61 62 3.49785 $w=1.3e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1005
+ $Y=0.2340 $X2=0.0855 $Y2=0.2340
r12 60 61 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1255
+ $Y=0.2340 $X2=0.1005 $Y2=0.2340
r13 15 22 3.36447 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1565 $Y=0.2340 $X2=0.1780 $Y2=0.2340
r14 15 60 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1565
+ $Y=0.2340 $X2=0.1255 $Y2=0.2340
r15 56 57 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r16 16 20 3.36447 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1565 $Y=0.0360 $X2=0.1780 $Y2=0.0360
r17 16 57 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1565
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r18 22 55 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.2340 $X2=0.1780 $Y2=0.2160
r19 20 52 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0360 $X2=0.1780 $Y2=0.0540
r20 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1980 $X2=0.1780 $Y2=0.2160
r21 53 54 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1865 $X2=0.1780 $Y2=0.1980
r22 18 21 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1780 $Y=0.1640 $X2=0.1780 $Y2=0.1350
r23 18 53 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1640 $X2=0.1780 $Y2=0.1865
r24 51 52 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0720 $X2=0.1780 $Y2=0.0540
r25 50 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.0835 $X2=0.1780 $Y2=0.0720
r26 17 21 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1780 $Y=0.1060 $X2=0.1780 $Y2=0.1350
r27 17 50 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1780
+ $Y=0.1060 $X2=0.1780 $Y2=0.0835
r28 12 41 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r29 9 35 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r30 44 45 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2055
+ $Y=0.1350 $X2=0.2145 $Y2=0.1350
r31 19 44 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1955
+ $Y=0.1350 $X2=0.2055 $Y2=0.1350
r32 19 21 2.90051 $w=1.55714e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1955 $Y=0.1350 $X2=0.1780 $Y2=0.1350
r33 10 28 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r34 39 41 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r35 38 39 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r36 37 38 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r37 33 35 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r38 31 32 7.08868 $w=1.53e-08 $l=1.2e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2130 $Y=0.1350 $X2=0.2250 $Y2=0.1350
r39 31 33 6.79332 $w=1.53e-08 $l=1.15e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2130 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r40 31 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2130 $Y=0.1350
+ $X2=0.2145 $Y2=0.1350
r41 29 32 3.24898 $w=1.53e-08 $l=5.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2250 $Y2=0.1350
r42 28 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r43 26 28 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2430 $Y2=0.1350
r44 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r45 24 25 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r46 11 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r47 1 24 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r48 1 37 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r49 11 24 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r50 11 37 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r51 3 14 1e-05
.ends

.subckt PM_OR2x4_ASAP7_75t_R%Y VSS 48 34 35 43 44 58 59 62 63 13 2 1 14 15 16
+ 17 27 26 3 4 18
c1 1 VSS 0.00846338f
c2 2 VSS 0.00845708f
c3 3 VSS 0.00849616f
c4 4 VSS 0.00851592f
c5 13 VSS 0.00454002f
c6 14 VSS 0.00443711f
c7 15 VSS 0.00451926f
c8 16 VSS 0.00442419f
c9 17 VSS 0.00127749f
c10 18 VSS 0.00107672f
c11 19 VSS 0.00906979f
c12 20 VSS 0.00911888f
c13 21 VSS 0.00108867f
c14 22 VSS 0.00109904f
c15 23 VSS 0.00648978f
c16 24 VSS 0.00648978f
c17 25 VSS 0.00731794f
c18 26 VSS 0.00233865f
c19 27 VSS 0.0026069f
c20 28 VSS 0.00218176f
c21 29 VSS 0.00218176f
c22 30 VSS 0.00345591f
c23 31 VSS 0.00345591f
r1 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 2 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 62 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 2 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 4 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r8 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r9 58 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r10 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1980 $X2=0.2160 $Y2=0.2160
r11 18 54 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1865 $X2=0.2160 $Y2=0.1980
r12 4 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.1980
r13 27 51 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2260 $Y2=0.2340
r14 27 55 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.2160 $Y2=0.2160
r15 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1980 $X2=0.3240 $Y2=0.2160
r16 22 52 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1865 $X2=0.3240 $Y2=0.1980
r17 20 29 11.1788 $w=1.38491e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2710 $Y=0.2340 $X2=0.3240 $Y2=0.2340
r18 20 51 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2710
+ $Y=0.2340 $X2=0.2260 $Y2=0.2340
r19 29 53 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3240 $Y2=0.2160
r20 24 31 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3645 $Y=0.2340 $X2=0.4050 $Y2=0.2340
r21 24 29 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3645 $Y=0.2340 $X2=0.3240 $Y2=0.2340
r22 31 50 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.4050 $Y2=0.2045
r23 49 50 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1660 $X2=0.4050 $Y2=0.2045
r24 48 49 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1475 $X2=0.4050 $Y2=0.1660
r25 48 47 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1475 $X2=0.4050 $Y2=0.1455
r26 46 47 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1455
r27 45 46 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1060 $X2=0.4050 $Y2=0.1350
r28 25 30 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0655 $X2=0.4050 $Y2=0.0360
r29 25 45 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0655 $X2=0.4050 $Y2=0.1060
r30 44 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r31 3 42 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r32 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r33 43 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r34 3 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0720
r35 23 28 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3645 $Y=0.0360 $X2=0.3240 $Y2=0.0360
r36 23 30 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3645 $Y=0.0360 $X2=0.4050 $Y2=0.0360
r37 21 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0540 $X2=0.3240 $Y2=0.0720
r38 21 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0540 $X2=0.3240 $Y2=0.0360
r39 28 38 11.1788 $w=1.38491e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.0360 $X2=0.2710 $Y2=0.0360
r40 19 26 0.682785 $w=1.75e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2260
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r41 19 38 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2260
+ $Y=0.0360 $X2=0.2710 $Y2=0.0360
r42 17 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0720
r43 17 26 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0360
r44 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0720
r45 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r46 1 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r47 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r48 34 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
.ends


*
.SUBCKT OR2x4_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 VSS N_MM5_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@4 VSS N_MM5@4_g N_MM5@4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 VSS N_MM0@3_g N_MM5@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 VSS N_MM0@2_g N_MM5@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM1_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM2_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VDD N_MM5_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@4 VDD N_MM5@4_g N_MM0@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 VDD N_MM0@3_g N_MM0@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 VDD N_MM0@2_g N_MM0@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR2x4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR2x4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR2x4_ASAP7_75t_R%NET15 VSS N_MM4_d N_MM3_s N_NET15_1
+ PM_OR2x4_ASAP7_75t_R%NET15
cc_1 N_NET15_1 N_MM1_g 0.0174089f
cc_2 N_NET15_1 N_MM2_g 0.0173663f
x_PM_OR2x4_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_OR2x4_ASAP7_75t_R%noxref_9
cc_3 N_noxref_9_1 N_MM1_g 0.00248547f
cc_4 N_noxref_9_1 N_NET7_14 0.0372583f
cc_5 N_noxref_9_1 N_noxref_8_1 0.00185614f
x_PM_OR2x4_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1 PM_OR2x4_ASAP7_75t_R%noxref_8
cc_6 N_noxref_8_1 N_MM1_g 0.004668f
cc_7 N_noxref_8_1 N_NET7_13 0.000590618f
x_PM_OR2x4_ASAP7_75t_R%A VSS A N_MM2_g N_A_1 N_A_5 N_A_6 PM_OR2x4_ASAP7_75t_R%A
cc_8 N_MM2_g N_B_6 0.000834962f
cc_9 N_A_1 N_B_1 0.00177232f
cc_10 N_A N_B_6 0.00180613f
cc_11 N_MM2_g N_MM1_g 0.00839362f
x_PM_OR2x4_ASAP7_75t_R%B VSS B N_MM1_g N_B_6 N_B_1 N_B_7 N_B_5
+ PM_OR2x4_ASAP7_75t_R%B
x_PM_OR2x4_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR2x4_ASAP7_75t_R%noxref_10
cc_12 N_noxref_10_1 N_MM0@2_g 0.00145614f
cc_13 N_noxref_10_1 N_Y_14 0.000831502f
x_PM_OR2x4_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR2x4_ASAP7_75t_R%noxref_11
cc_14 N_noxref_11_1 N_MM0@2_g 0.00146161f
cc_15 N_noxref_11_1 N_Y_16 0.000831917f
cc_16 N_noxref_11_1 N_noxref_10_1 0.00178873f
x_PM_OR2x4_ASAP7_75t_R%NET7 VSS N_MM5_g N_MM5@4_g N_MM0@3_g N_MM0@2_g N_MM1_s
+ N_MM2_s N_MM4_s N_NET7_13 N_NET7_16 N_NET7_3 N_NET7_4 N_NET7_15 N_NET7_14
+ N_NET7_1 N_NET7_21 N_NET7_17 N_NET7_18 N_NET7_22 N_NET7_20 N_NET7_19
+ PM_OR2x4_ASAP7_75t_R%NET7
cc_17 N_NET7_13 N_MM1_g 0.0113412f
cc_18 N_NET7_16 N_MM1_g 0.000387338f
cc_19 N_NET7_3 N_B_6 0.000420777f
cc_20 N_NET7_3 N_B_1 0.000533292f
cc_21 N_NET7_4 N_MM1_g 0.000609965f
cc_22 N_NET7_16 N_B_7 0.000830889f
cc_23 N_NET7_15 N_B_5 0.000962122f
cc_24 N_NET7_3 N_B_5 0.00162267f
cc_25 N_NET7_14 N_B_1 0.00195472f
cc_26 N_NET7_3 N_MM1_g 0.00250821f
cc_27 N_NET7_14 N_MM1_g 0.0502572f
cc_28 N_NET7_13 N_MM2_g 0.0114005f
cc_29 N_NET7_3 N_MM2_g 0.000410267f
cc_30 N_NET7_1 N_MM2_g 0.000431869f
cc_31 N_NET7_21 N_MM2_g 0.000571122f
cc_32 N_NET7_1 N_A_1 0.000773389f
cc_33 N_NET7_4 N_MM2_g 0.00080444f
cc_34 N_NET7_17 N_A 0.00188632f
cc_35 N_NET7_18 N_A 0.00202415f
cc_36 N_NET7_21 N_A 0.00450556f
cc_37 N_NET7_16 N_A_5 0.00499563f
cc_38 N_NET7_15 N_A_6 0.00500908f
cc_39 N_MM5_g N_MM2_g 0.018002f
x_PM_OR2x4_ASAP7_75t_R%Y VSS Y N_MM5_s N_MM5@4_s N_MM5@3_s N_MM5@2_s N_MM0@3_s
+ N_MM0@2_s N_MM0_s N_MM0@4_s N_Y_13 N_Y_2 N_Y_1 N_Y_14 N_Y_15 N_Y_16 N_Y_17
+ N_Y_27 N_Y_26 N_Y_3 N_Y_4 N_Y_18 PM_OR2x4_ASAP7_75t_R%Y
cc_40 N_Y_13 N_NET7_1 0.00105385f
cc_41 N_Y_13 N_NET7_22 0.000295477f
cc_42 N_Y_13 N_NET7_20 0.000303371f
cc_43 N_Y_2 N_NET7_18 0.00063231f
cc_44 N_Y_1 N_NET7_17 0.000643327f
cc_45 N_Y_14 N_MM0@2_g 0.0676843f
cc_46 N_Y_15 N_MM5@4_g 0.0308014f
cc_47 N_Y_16 N_MM0@2_g 0.0308163f
cc_48 N_Y_1 N_NET7_1 0.000923611f
cc_49 N_Y_17 N_NET7_19 0.0011842f
cc_50 N_Y_27 N_NET7_22 0.001627f
cc_51 N_Y_26 N_NET7_20 0.00165363f
cc_52 N_Y_3 N_MM0@2_g 0.00174613f
cc_53 N_Y_4 N_MM0@2_g 0.0017517f
cc_54 N_Y_2 N_MM5@4_g 0.00214179f
cc_55 N_Y_1 N_MM5@4_g 0.00223283f
cc_56 N_Y_17 N_NET7_17 0.00411628f
cc_57 N_Y_18 N_NET7_18 0.00412911f
cc_58 N_Y_16 N_NET7_1 0.00958589f
cc_59 N_Y_13 N_MM5_g 0.0368878f
cc_60 N_Y_14 N_MM0@3_g 0.036975f
cc_61 N_Y_13 N_MM5@4_g 0.0687984f
*END of OR2x4_ASAP7_75t_R.pxi
.ENDS
** Design:	OR2x6_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR2x6_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR2x6_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR2x6_ASAP7_75t_R%NET15 VSS 2 3 1
c1 1 VSS 0.000944831f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_OR2x6_ASAP7_75t_R%noxref_9 VSS 1
c1 1 VSS 0.0323233f
.ends

.subckt PM_OR2x6_ASAP7_75t_R%NET15__2 VSS 2 3 1
c1 1 VSS 0.000908052f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR2x6_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0421287f
.ends

.subckt PM_OR2x6_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0423141f
.ends

.subckt PM_OR2x6_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0423578f
.ends

.subckt PM_OR2x6_ASAP7_75t_R%Y VSS 40 32 33 44 45 48 49 60 61 64 65 68 69 19 27
+ 26 25 21 20 22 24 23 2 5 6 4 3 1
c1 1 VSS 0.0101797f
c2 2 VSS 0.00984167f
c3 3 VSS 0.00989334f
c4 4 VSS 0.0102651f
c5 5 VSS 0.00984703f
c6 6 VSS 0.00979525f
c7 19 VSS 0.00450362f
c8 20 VSS 0.00438423f
c9 21 VSS 0.00440818f
c10 22 VSS 0.0044351f
c11 23 VSS 0.00440505f
c12 24 VSS 0.00442128f
c13 25 VSS 0.0317792f
c14 26 VSS 0.0297806f
c15 27 VSS 0.00747662f
c16 28 VSS 0.00336908f
c17 29 VSS 0.00333577f
r1 69 67 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r2 6 67 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r3 24 6 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r4 68 24 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
r5 65 63 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 4 63 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 23 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 64 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r10 2 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r11 22 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r12 60 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r13 6 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5400 $Y2=0.2340
r14 4 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r15 2 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r16 54 55 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.2340 $X2=0.5805 $Y2=0.2340
r17 53 54 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5400 $Y2=0.2340
r18 52 53 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r19 51 52 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r20 50 51 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r21 25 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r22 29 41 9.4274 $w=1.48568e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.6210 $Y2=0.1865
r23 29 55 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.2340 $X2=0.5805 $Y2=0.2340
r24 49 47 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r25 5 47 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r26 21 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r27 48 21 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r28 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r29 3 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r30 20 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r31 44 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r32 40 41 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1475 $X2=0.6210 $Y2=0.1865
r33 40 27 12.0093 $w=1.3e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1475 $X2=0.6210 $Y2=0.0960
r34 27 28 12.3423 $w=1.447e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0960 $X2=0.6210 $Y2=0.0360
r35 5 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5400 $Y2=0.0360
r36 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r37 28 39 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.0360 $X2=0.5805 $Y2=0.0360
r38 38 39 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5400
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r39 37 38 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5400 $Y2=0.0360
r40 36 37 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r41 35 36 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r42 34 35 12.5922 $w=1.3e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r43 26 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3125
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r44 1 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r45 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r46 1 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r47 19 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r48 32 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
.ends

.subckt PM_OR2x6_ASAP7_75t_R%A VSS 32 3 4 5 6 7 1 9
c1 1 VSS 0.00526106f
c2 3 VSS 0.0322904f
c3 4 VSS 0.0324257f
c4 5 VSS 0.0211851f
c5 6 VSS 0.00555889f
c6 7 VSS 0.00169685f
c7 8 VSS 0.00407449f
c8 9 VSS 0.000518281f
r1 32 31 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1340 $X2=0.0270 $Y2=0.1197
r2 5 8 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0935 $X2=0.0270 $Y2=0.0720
r3 5 31 6.12123 $w=1.3e-08 $l=2.62e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0935 $X2=0.0270 $Y2=0.1197
r4 8 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0720 $X2=0.0540 $Y2=0.0720
r5 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0540 $Y2=0.0720
r6 28 29 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0920
+ $Y=0.0720 $X2=0.0810 $Y2=0.0720
r7 6 9 4.29228 $w=1.42791e-08 $l=2.52438e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1100 $Y=0.0720 $X2=0.1350 $Y2=0.0755
r8 6 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1100
+ $Y=0.0720 $X2=0.0920 $Y2=0.0720
r9 9 22 1.37741 $w=1.60556e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0755 $X2=0.1350 $Y2=0.0845
r10 4 19 2.92627 $w=1.245e-07 $l=2.7e-08 $layer=LIG $thickness=5.2e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1080
r11 21 23 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1025 $X2=0.1350 $Y2=0.1115
r12 7 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0935 $X2=0.1350 $Y2=0.1025
r13 7 22 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0935 $X2=0.1350 $Y2=0.0845
r14 17 19 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1080 $X2=0.1890 $Y2=0.1080
r15 16 17 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1080 $X2=0.1765 $Y2=0.1080
r16 15 16 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1080 $X2=0.1620 $Y2=0.1080
r17 13 15 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1445 $Y=0.1080 $X2=0.1475 $Y2=0.1080
r18 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1080 $X2=0.1445 $Y2=0.1080
r19 12 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1080
+ $X2=0.1350 $Y2=0.1115
r20 1 12 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1080 $X2=0.1350 $Y2=0.1080
r21 1 14 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1080 $X2=0.1245 $Y2=0.1080
r22 11 12 2.35044 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1080 $X2=0.1350 $Y2=0.1080
r23 11 14 0.295362 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1080 $X2=0.1245 $Y2=0.1080
r24 11 15 1.47681 $w=1.53e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1350 $Y=0.1080 $X2=0.1475 $Y2=0.1080
r25 3 11 0.314665 $w=2.27e-07 $l=2.7e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1080
.ends

.subckt PM_OR2x6_ASAP7_75t_R%B VSS 22 5 6 1 8 7 9 10 11 2
c1 1 VSS 0.00465568f
c2 2 VSS 0.00597588f
c3 5 VSS 0.0720639f
c4 6 VSS 0.0826806f
c5 7 VSS 0.00149567f
c6 8 VSS 0.00590131f
c7 9 VSS 0.00253167f
c8 10 VSS 0.00120993f
c9 11 VSS 0.0020348f
r1 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1485
r4 11 23 8.08899 $w=1.41321e-08 $l=3.98e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1620 $X2=0.2032 $Y2=0.1620
r5 11 26 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1620 $X2=0.2430 $Y2=0.1485
r6 22 23 7.28718 $w=1.3e-08 $l=3.12e-08 $layer=M1 $thickness=3.6e-08 $X=0.1720
+ $Y=0.1620 $X2=0.2032 $Y2=0.1620
r7 22 21 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.1720
+ $Y=0.1620 $X2=0.1597 $Y2=0.1620
r8 20 21 3.20636 $w=1.3e-08 $l=1.37e-08 $layer=M1 $thickness=3.6e-08 $X=0.1460
+ $Y=0.1620 $X2=0.1597 $Y2=0.1620
r9 19 20 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1620 $X2=0.1460 $Y2=0.1620
r10 9 10 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.1620 $X2=0.0810 $Y2=0.1620
r11 9 19 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1620 $X2=0.1350 $Y2=0.1620
r12 8 10 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1800 $X2=0.0810 $Y2=0.1620
r13 10 15 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1620 $X2=0.0810 $Y2=0.1485
r14 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1485
r15 13 14 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1240 $X2=0.0810 $Y2=0.1350
r16 7 13 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1140 $X2=0.0810 $Y2=0.1240
r17 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r18 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_OR2x6_ASAP7_75t_R%NET7 VSS 12 13 14 15 16 17 81 82 90 91 94 95 20 24
+ 19 1 5 22 3 27 4 25 18 21 28 29
c1 1 VSS 0.030324f
c2 3 VSS 0.011507f
c3 4 VSS 0.00840817f
c4 5 VSS 0.011384f
c5 12 VSS 0.0820011f
c6 13 VSS 0.0818314f
c7 14 VSS 0.081777f
c8 15 VSS 0.0817465f
c9 16 VSS 0.0816184f
c10 17 VSS 0.082316f
c11 18 VSS 0.00840649f
c12 19 VSS 0.0084175f
c13 20 VSS 0.00745684f
c14 21 VSS 0.0149643f
c15 22 VSS 0.00773564f
c16 23 VSS 0.00236468f
c17 24 VSS 0.00284158f
c18 25 VSS 0.00369285f
c19 26 VSS 0.00430713f
c20 27 VSS 0.00204353f
c21 28 VSS 0.00216857f
c22 29 VSS 0.00214805f
r1 95 93 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r2 3 93 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r3 18 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r4 94 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r5 91 89 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r6 5 89 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0540 $X2=0.2305 $Y2=0.0540
r7 19 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0540 $X2=0.2160 $Y2=0.0540
r8 90 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0540 $X2=0.2015 $Y2=0.0540
r9 3 86 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1080 $Y2=0.0360
r10 5 83 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r11 86 87 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r12 83 84 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r13 21 83 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r14 21 87 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r15 26 78 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2430 $Y2=0.0540
r16 26 84 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0360 $X2=0.2295 $Y2=0.0360
r17 82 80 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r18 4 80 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.2025 $X2=0.1765 $Y2=0.2025
r19 20 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r20 81 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r21 23 27 1.37741 $w=1.60556e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0665 $X2=0.2430 $Y2=0.0755
r22 23 78 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0665 $X2=0.2430 $Y2=0.0540
r23 4 75 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.2025
+ $X2=0.1620 $Y2=0.1980
r24 75 76 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.1980 $X2=0.2025 $Y2=0.1980
r25 73 76 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2025 $Y2=0.1980
r26 22 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1980 $X2=0.2970 $Y2=0.1980
r27 22 73 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r28 24 28 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.0790 $X2=0.2970 $Y2=0.0790
r29 24 27 4.75866 $w=1.41702e-08 $l=2.72259e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.0790 $X2=0.2430 $Y2=0.0755
r30 29 67 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2970 $Y2=0.1800
r31 17 62 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r32 16 56 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r33 15 50 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r34 14 44 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r35 13 38 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r36 66 67 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1575 $X2=0.2970 $Y2=0.1800
r37 65 66 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1575
r38 64 65 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1235 $X2=0.2970 $Y2=0.1350
r39 25 64 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1045 $X2=0.2970 $Y2=0.1235
r40 25 28 4.29723 $w=1.64588e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1045 $X2=0.2970 $Y2=0.0790
r41 60 62 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5545 $Y=0.1350 $X2=0.5670 $Y2=0.1350
r42 59 60 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5400 $Y=0.1350 $X2=0.5545 $Y2=0.1350
r43 57 59 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5255 $Y=0.1350 $X2=0.5400 $Y2=0.1350
r44 56 57 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5130 $Y=0.1350 $X2=0.5255 $Y2=0.1350
r45 54 56 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r46 53 54 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r47 51 53 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r48 50 51 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r49 48 50 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r50 47 48 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r51 45 47 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r52 44 45 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r53 42 44 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r54 41 42 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r55 39 41 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r56 38 39 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r57 36 38 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r58 35 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r59 34 35 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r60 32 34 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r61 31 32 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r62 31 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
r63 1 31 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r64 1 33 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2865 $Y2=0.1350
r65 12 31 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r66 12 33 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2970 $Y=0.1350 $X2=0.2865 $Y2=0.1350
r67 12 34 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
.ends


*
.SUBCKT OR2x6_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 VSS N_MM4@2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2@2 VSS N_MM4_g N_MM2@2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1@2 VSS N_MM3_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM5 VSS N_MM0_g N_MM5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@6 VSS N_MM0@6_g N_MM5@6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@5 VSS N_MM0@5_g N_MM5@5_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@4 VSS N_MM0@4_g N_MM5@4_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@3 VSS N_MM0@3_g N_MM5@3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 VSS N_MM0@2_g N_MM5@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3@2 VDD N_MM1_g N_MM3@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 VDD N_MM0_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@6 VDD N_MM0@6_g N_MM0@6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@5 VDD N_MM0@5_g N_MM0@5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@4 VDD N_MM0@4_g N_MM0@4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 VDD N_MM0@3_g N_MM0@3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 VDD N_MM0@2_g N_MM0@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR2x6_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR2x6_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR2x6_ASAP7_75t_R%NET15 VSS N_MM4_d N_MM3_s N_NET15_1
+ PM_OR2x6_ASAP7_75t_R%NET15
cc_1 N_NET15_1 N_MM3_g 0.0174337f
cc_2 N_NET15_1 N_MM4_g 0.0173723f
x_PM_OR2x6_ASAP7_75t_R%noxref_9 VSS N_noxref_9_1 PM_OR2x6_ASAP7_75t_R%noxref_9
cc_3 N_noxref_9_1 N_MM1_g 0.00346687f
cc_4 N_noxref_9_1 N_MM4@2_g 0.000897109f
x_PM_OR2x6_ASAP7_75t_R%NET15__2 VSS N_MM3@2_s N_MM4@2_d N_NET15__2_1
+ PM_OR2x6_ASAP7_75t_R%NET15__2
cc_5 N_NET15__2_1 N_MM1_g 0.0171643f
cc_6 N_NET15__2_1 N_MM4@2_g 0.0172408f
x_PM_OR2x6_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR2x6_ASAP7_75t_R%noxref_10
cc_7 N_noxref_10_1 N_MM1_g 0.00161168f
cc_8 N_noxref_10_1 N_MM4@2_g 0.000803006f
cc_9 N_noxref_10_1 N_noxref_9_1 0.00189333f
x_PM_OR2x6_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR2x6_ASAP7_75t_R%noxref_11
cc_10 N_noxref_11_1 N_MM0@2_g 0.00145309f
cc_11 N_noxref_11_1 N_Y_21 0.00083652f
x_PM_OR2x6_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR2x6_ASAP7_75t_R%noxref_12
cc_12 N_noxref_12_1 N_MM0@2_g 0.00146199f
cc_13 N_noxref_12_1 N_Y_24 0.000849847f
cc_14 N_noxref_12_1 N_noxref_11_1 0.0017765f
x_PM_OR2x6_ASAP7_75t_R%Y VSS Y N_MM5_s N_MM5@6_s N_MM5@5_s N_MM5@4_s N_MM5@3_s
+ N_MM5@2_s N_MM0_s N_MM0@6_s N_MM0@5_s N_MM0@4_s N_MM0@3_s N_MM0@2_s N_Y_19
+ N_Y_27 N_Y_26 N_Y_25 N_Y_21 N_Y_20 N_Y_22 N_Y_24 N_Y_23 N_Y_2 N_Y_5 N_Y_6
+ N_Y_4 N_Y_3 N_Y_1 PM_OR2x6_ASAP7_75t_R%Y
cc_15 N_Y_19 N_NET7_24 0.000282775f
cc_16 N_Y_19 N_NET7_1 0.00040452f
cc_17 N_Y_27 N_NET7_1 0.000515816f
cc_18 N_Y_26 N_NET7_28 0.00072885f
cc_19 N_Y_25 N_NET7_22 0.000775406f
cc_20 N_Y_21 N_MM0@2_g 0.0669953f
cc_21 N_Y_20 N_MM0@4_g 0.0671775f
cc_22 N_Y_22 N_MM0@6_g 0.0304842f
cc_23 N_Y_24 N_MM0@2_g 0.0303901f
cc_24 N_Y_23 N_MM0@4_g 0.0305797f
cc_25 N_Y_25 N_NET7_29 0.00129096f
cc_26 N_Y_2 N_NET7_25 0.0014319f
cc_27 N_Y_26 N_MM0@4_g 0.0016581f
cc_28 N_Y_5 N_MM0@2_g 0.00180697f
cc_29 N_Y_6 N_MM0@2_g 0.00181144f
cc_30 N_Y_4 N_MM0@4_g 0.00186672f
cc_31 N_Y_3 N_MM0@4_g 0.0018856f
cc_32 N_Y_2 N_MM0@6_g 0.00233986f
cc_33 N_Y_1 N_MM0@6_g 0.00236204f
cc_34 N_Y_25 N_MM0@4_g 0.00239628f
cc_35 N_Y_23 N_NET7_1 0.0149977f
cc_36 N_Y_19 N_MM0_g 0.0365477f
cc_37 N_Y_21 N_MM0@3_g 0.0366444f
cc_38 N_Y_20 N_MM0@5_g 0.0366581f
cc_39 N_Y_19 N_MM0@6_g 0.0683265f
x_PM_OR2x6_ASAP7_75t_R%A VSS A N_MM4@2_g N_MM4_g N_A_5 N_A_6 N_A_7 N_A_1 N_A_9
+ PM_OR2x6_ASAP7_75t_R%A
cc_40 N_A_5 N_MM1_g 0.000790114f
cc_41 N_MM4@2_g N_B_1 0.000816019f
cc_42 N_A_5 N_B_8 0.00123798f
cc_43 N_A_6 N_B_7 0.00128196f
cc_44 N_A_7 N_B_7 0.00155936f
cc_45 N_A_1 N_MM3_g 0.00177221f
cc_46 N_A_7 N_B_9 0.00197508f
cc_47 N_A_5 N_B_7 0.00249143f
cc_48 N_A_5 N_B_10 0.00348136f
cc_49 N_MM4_g N_MM3_g 0.00720284f
cc_50 N_MM4@2_g N_MM1_g 0.00913367f
x_PM_OR2x6_ASAP7_75t_R%B VSS B N_MM1_g N_MM3_g N_B_1 N_B_8 N_B_7 N_B_9 N_B_10
+ N_B_11 N_B_2 PM_OR2x6_ASAP7_75t_R%B
x_PM_OR2x6_ASAP7_75t_R%NET7 VSS N_MM0_g N_MM0@6_g N_MM0@5_g N_MM0@4_g N_MM0@3_g
+ N_MM0@2_g N_MM4@2_s N_MM4_s N_MM2@2_s N_MM1@2_s N_MM1_s N_MM2_s N_NET7_20
+ N_NET7_24 N_NET7_19 N_NET7_1 N_NET7_5 N_NET7_22 N_NET7_3 N_NET7_27 N_NET7_4
+ N_NET7_25 N_NET7_18 N_NET7_21 N_NET7_28 N_NET7_29 PM_OR2x6_ASAP7_75t_R%NET7
cc_51 N_NET7_20 N_MM1_g 0.000304873f
cc_52 N_NET7_24 N_MM1_g 0.000334321f
cc_53 N_NET7_19 N_MM1_g 0.000351062f
cc_54 N_NET7_1 N_MM3_g 0.000433958f
cc_55 N_NET7_5 N_MM3_g 0.00047166f
cc_56 N_NET7_22 N_B_8 0.000475171f
cc_57 N_NET7_3 N_MM1_g 0.000476402f
cc_58 N_NET7_27 N_B_11 0.000538185f
cc_59 N_NET7_4 N_B_9 0.00185033f
cc_60 N_NET7_1 N_B_2 0.00201427f
cc_61 N_NET7_22 N_B_11 0.00111297f
cc_62 N_NET7_25 N_B_11 0.00278921f
cc_63 N_NET7_19 N_MM3_g 0.0109725f
cc_64 N_NET7_22 N_B_9 0.00989324f
cc_65 N_MM0_g N_MM3_g 0.0172428f
cc_66 N_NET7_18 N_MM1_g 0.0262983f
cc_67 N_NET7_19 N_MM4_g 0.0114497f
cc_68 N_NET7_18 N_MM4_g 0.00035906f
cc_69 N_NET7_3 N_MM4_g 0.000411824f
cc_70 N_NET7_3 N_A_6 0.000432635f
cc_71 N_NET7_21 N_A_7 0.000567323f
cc_72 N_NET7_5 N_MM4_g 0.000837686f
cc_73 N_NET7_3 N_MM4@2_g 0.00136656f
cc_74 N_NET7_4 N_MM4_g 0.00148919f
cc_75 N_NET7_21 N_A_6 0.00233884f
cc_76 N_NET7_19 N_A_1 0.00269486f
cc_77 N_NET7_18 N_MM4@2_g 0.011119f
cc_78 N_NET7_21 N_A_9 0.00417488f
cc_79 N_NET7_20 N_MM4@2_g 0.0332049f
cc_80 N_NET7_20 N_MM4_g 0.0660341f
*END of OR2x6_ASAP7_75t_R.pxi
.ENDS
** Design:	OR3x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR3x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR3x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR3x1_ASAP7_75t_R%NET67 VSS 2 3 1
c1 1 VSS 0.000975174f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR3x1_ASAP7_75t_R%NET66 VSS 2 3 1
c1 1 VSS 0.000966236f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR3x1_ASAP7_75t_R%B VSS 6 3 1 4
c1 1 VSS 0.00599243f
c2 3 VSS 0.0461347f
c3 4 VSS 0.00424848f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_OR3x1_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00476142f
.ends

.subckt PM_OR3x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00502891f
.ends

.subckt PM_OR3x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00486012f
.ends

.subckt PM_OR3x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00471181f
.ends

.subckt PM_OR3x1_ASAP7_75t_R%C VSS 4 3 1
c1 1 VSS 0.00622298f
c2 3 VSS 0.0830003f
c3 4 VSS 0.00418069f
r1 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 4 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_OR3x1_ASAP7_75t_R%A VSS 6 3 1 4
c1 1 VSS 0.00265841f
c2 3 VSS 0.0429958f
c3 4 VSS 0.0121946f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1355
.ends

.subckt PM_OR3x1_ASAP7_75t_R%Y VSS 23 15 30 7 9 1 2 8 11 10 12
c1 1 VSS 0.00688839f
c2 2 VSS 0.00727915f
c3 7 VSS 0.00365809f
c4 8 VSS 0.00360518f
c5 9 VSS 0.00297253f
c6 10 VSS 0.00131001f
c7 11 VSS 0.00157104f
c8 12 VSS 0.00269083f
c9 13 VSS 0.000888302f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2680 $Y2=0.2025
r2 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r3 2 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2170
r4 26 27 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2045 $X2=0.2700 $Y2=0.2170
r5 12 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.1920 $X2=0.2835 $Y2=0.1920
r6 12 26 1.73456 $w=1.66e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1920 $X2=0.2700 $Y2=0.2045
r7 13 24 4.99922 $w=1.46981e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1920 $X2=0.2970 $Y2=0.1655
r8 13 25 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1920 $X2=0.2835 $Y2=0.1920
r9 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1655
r10 23 22 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1475 $X2=0.2970 $Y2=0.1455
r11 21 22 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1455
r12 10 20 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1100 $X2=0.2970 $Y2=0.0850
r13 10 21 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1100 $X2=0.2970 $Y2=0.1350
r14 19 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2835 $Y=0.0850 $X2=0.2970 $Y2=0.0850
r15 18 19 1.91673 $w=1.62692e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2705 $Y=0.0850 $X2=0.2835 $Y2=0.0850
r16 11 17 0.867186 $w=1.3625e-08 $l=1.51162e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2615 $Y=0.0850 $X2=0.2700 $Y2=0.0725
r17 11 18 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2615
+ $Y=0.0850 $X2=0.2705 $Y2=0.0850
r18 16 17 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0600 $X2=0.2700 $Y2=0.0725
r19 9 16 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0425 $X2=0.2700 $Y2=0.0600
r20 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0600
r21 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2680 $Y2=0.0675
r22 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_OR3x1_ASAP7_75t_R%NET61 VSS 12 60 61 63 65 15 3 16 17 4 13 5 14 1 21
+ 18 19 22 20
c1 1 VSS 0.00358393f
c2 3 VSS 0.00861801f
c3 4 VSS 0.00642461f
c4 5 VSS 0.00983709f
c5 12 VSS 0.0804683f
c6 13 VSS 0.00401072f
c7 14 VSS 0.0050046f
c8 15 VSS 0.0030881f
c9 16 VSS 0.0169715f
c10 17 VSS 0.0178347f
c11 18 VSS 0.00213392f
c12 19 VSS 0.00221967f
c13 20 VSS 0.00271258f
c14 21 VSS 0.000398974f
c15 22 VSS 0.00315028f
r1 65 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 15 64 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 63 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r4 13 62 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r5 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 5 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 14 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 60 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r10 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r11 5 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r12 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 54 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 51 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 17 22 2.60893 $w=1.47857e-08 $l=1.84391e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2070 $Y=0.2340 $X2=0.2250 $Y2=0.2300
r19 17 50 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r20 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r21 46 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r22 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r23 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r24 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r25 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r26 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r27 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r28 16 20 2.65995 $w=1.48966e-08 $l=1.83371e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2070 $Y=0.0360 $X2=0.2250 $Y2=0.0395
r29 16 40 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2070
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 22 37 3.42509 $w=1.44286e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.2300 $X2=0.2250 $Y2=0.2125
r31 20 35 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.0395 $X2=0.2250 $Y2=0.0575
r32 36 37 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1915 $X2=0.2250 $Y2=0.2125
r33 19 21 5.4656 $w=1.45789e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1635 $X2=0.2250 $Y2=0.1350
r34 19 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1635 $X2=0.2250 $Y2=0.1915
r35 34 35 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0730 $X2=0.2250 $Y2=0.0575
r36 33 34 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.0850 $X2=0.2250 $Y2=0.0730
r37 18 21 4.64944 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1100 $X2=0.2250 $Y2=0.1350
r38 18 33 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2250
+ $Y=0.1100 $X2=0.2250 $Y2=0.0850
r39 29 30 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2365
+ $Y=0.1350 $X2=0.2480 $Y2=0.1350
r40 21 29 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2250 $Y=0.1350 $X2=0.2365 $Y2=0.1350
r41 24 26 3.00957 $w=2.05111e-08 $l=9e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2460 $Y=0.1350 $X2=0.2550 $Y2=0.1350
r42 24 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2460 $Y=0.1350
+ $X2=0.2480 $Y2=0.1350
r43 1 24 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2360
+ $Y=0.1350 $X2=0.2460 $Y2=0.1350
r44 1 25 1.07884 $w=2.10429e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2360 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r45 12 24 2.14279 $w=1.42588e-07 $l=3e-09 $layer=LIG $thickness=5.27059e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2460 $Y2=0.1350
r46 12 25 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r47 12 26 1.49611 $w=1.91717e-07 $l=1.2e-08 $layer=LIG $thickness=5.46667e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2550 $Y2=0.1350
r48 4 15 1e-05
r49 3 13 1e-05
.ends


*
.SUBCKT OR3x1_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM12_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR3x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR3x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR3x1_ASAP7_75t_R%NET67 VSS N_MM11_s N_MM10_d N_NET67_1
+ PM_OR3x1_ASAP7_75t_R%NET67
cc_1 N_NET67_1 N_MM12_g 0.0172626f
cc_2 N_NET67_1 N_MM13_g 0.0172437f
x_PM_OR3x1_ASAP7_75t_R%NET66 VSS N_MM10_s N_MM8_d N_NET66_1
+ PM_OR3x1_ASAP7_75t_R%NET66
cc_3 N_NET66_1 N_MM13_g 0.0173629f
cc_4 N_NET66_1 N_MM14_g 0.0172334f
x_PM_OR3x1_ASAP7_75t_R%B VSS B N_MM13_g N_B_1 N_B_4 PM_OR3x1_ASAP7_75t_R%B
cc_5 N_B_1 N_A_1 0.00131253f
cc_6 N_B_4 N_A_4 0.00472198f
cc_7 N_MM13_g N_MM12_g 0.00609968f
x_PM_OR3x1_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR3x1_ASAP7_75t_R%noxref_10
cc_8 N_noxref_10_1 N_MM12_g 0.0016326f
cc_9 N_noxref_10_1 N_NET61_13 0.0381688f
x_PM_OR3x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR3x1_ASAP7_75t_R%noxref_11
cc_10 N_noxref_11_1 N_MM12_g 0.00163702f
cc_11 N_noxref_11_1 N_NET61_15 0.0378946f
cc_12 N_noxref_11_1 N_noxref_10_1 0.00179434f
x_PM_OR3x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_OR3x1_ASAP7_75t_R%noxref_13
cc_13 N_noxref_13_1 N_MM1_g 0.00148924f
cc_14 N_noxref_13_1 N_Y_8 0.0382988f
cc_15 N_noxref_13_1 N_noxref_12_1 0.00177898f
x_PM_OR3x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR3x1_ASAP7_75t_R%noxref_12
cc_16 N_noxref_12_1 N_MM1_g 0.00148261f
cc_17 N_noxref_12_1 N_Y_7 0.0383693f
x_PM_OR3x1_ASAP7_75t_R%C VSS C N_MM14_g N_C_1 PM_OR3x1_ASAP7_75t_R%C
cc_18 N_MM14_g N_B_1 0.00131113f
cc_19 N_C N_B_4 0.00488458f
cc_20 N_MM14_g N_MM13_g 0.00619531f
x_PM_OR3x1_ASAP7_75t_R%A VSS A N_MM12_g N_A_1 N_A_4 PM_OR3x1_ASAP7_75t_R%A
x_PM_OR3x1_ASAP7_75t_R%Y VSS Y N_MM1_d N_MM0_d N_Y_7 N_Y_9 N_Y_1 N_Y_2 N_Y_8
+ N_Y_11 N_Y_10 N_Y_12 PM_OR3x1_ASAP7_75t_R%Y
cc_21 N_Y_7 N_NET61_19 0.000380381f
cc_22 N_Y_7 N_NET61_18 0.000380478f
cc_23 N_Y_7 N_NET61_22 0.000511579f
cc_24 N_Y_9 N_NET61_20 0.000601772f
cc_25 N_Y_9 N_NET61_18 0.00110017f
cc_26 N_Y_1 N_NET61_1 0.00117971f
cc_27 N_Y_1 N_MM1_g 0.00133958f
cc_28 N_Y_2 N_MM1_g 0.00137464f
cc_29 N_Y_8 N_NET61_1 0.00219456f
cc_30 N_Y_11 N_NET61_18 0.0027628f
cc_31 N_Y_10 N_NET61_21 0.00294185f
cc_32 N_Y_12 N_NET61_19 0.00350625f
cc_33 N_Y_8 N_MM1_g 0.0151977f
cc_34 N_Y_7 N_MM1_g 0.0552148f
x_PM_OR3x1_ASAP7_75t_R%NET61 VSS N_MM1_g N_MM13_d N_MM14_d N_MM12_d N_MM11_d
+ N_NET61_15 N_NET61_3 N_NET61_16 N_NET61_17 N_NET61_4 N_NET61_13 N_NET61_5
+ N_NET61_14 N_NET61_1 N_NET61_21 N_NET61_18 N_NET61_19 N_NET61_22 N_NET61_20
+ PM_OR3x1_ASAP7_75t_R%NET61
cc_35 N_NET61_15 N_MM12_g 0.0158722f
cc_36 N_NET61_3 N_A_1 0.000634359f
cc_37 N_NET61_16 N_A_4 0.00130074f
cc_38 N_NET61_17 N_A_4 0.00139411f
cc_39 N_NET61_3 N_MM12_g 0.00154794f
cc_40 N_NET61_15 N_A_1 0.0016759f
cc_41 N_NET61_4 N_MM12_g 0.00188998f
cc_42 N_NET61_3 N_A_4 0.0042347f
cc_43 N_NET61_13 N_MM12_g 0.0549175f
cc_44 N_NET61_5 N_MM13_g 0.00152725f
cc_45 N_NET61_14 N_B_1 0.000915317f
cc_46 N_NET61_16 N_B_4 0.00119104f
cc_47 N_NET61_17 N_B_4 0.00144368f
cc_48 N_NET61_5 N_B_4 0.0033059f
cc_49 N_NET61_14 N_MM13_g 0.0360851f
cc_50 N_NET61_1 N_MM14_g 0.000464228f
cc_51 N_NET61_21 N_MM14_g 0.00081478f
cc_52 N_NET61_16 N_C 0.000909888f
cc_53 N_NET61_17 N_C 0.0010523f
cc_54 N_NET61_14 N_C_1 0.0011601f
cc_55 N_NET61_5 N_MM14_g 0.00119629f
cc_56 N_MM1_g N_MM14_g 0.00164215f
cc_57 N_NET61_18 N_C 0.00221207f
cc_58 N_NET61_19 N_C 0.00243677f
cc_59 N_NET61_21 N_C 0.00771242f
cc_60 N_NET61_14 N_MM14_g 0.0367682f
*END of OR3x1_ASAP7_75t_R.pxi
.ENDS
** Design:	OR3x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR3x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR3x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR3x2_ASAP7_75t_R%NET67 VSS 2 3 1
c1 1 VSS 0.000977234f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR3x2_ASAP7_75t_R%NET66 VSS 2 3 1
c1 1 VSS 0.000960302f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR3x2_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00480312f
.ends

.subckt PM_OR3x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0422942f
.ends

.subckt PM_OR3x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0422977f
.ends

.subckt PM_OR3x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00491486f
.ends

.subckt PM_OR3x2_ASAP7_75t_R%C VSS 7 3 4 1
c1 1 VSS 0.00673831f
c2 3 VSS 0.0830905f
c3 4 VSS 0.00454911f
r1 7 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 7 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_OR3x2_ASAP7_75t_R%A VSS 6 3 1 4
c1 1 VSS 0.00267877f
c2 3 VSS 0.0429845f
c3 4 VSS 0.0123838f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1355
.ends

.subckt PM_OR3x2_ASAP7_75t_R%B VSS 6 3 1 4
c1 1 VSS 0.00526928f
c2 3 VSS 0.0459214f
c3 4 VSS 0.00395527f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_OR3x2_ASAP7_75t_R%Y VSS 28 20 21 36 37 7 1 13 15 14 9 2 10 8
c1 1 VSS 0.00845752f
c2 2 VSS 0.00837598f
c3 7 VSS 0.0045721f
c4 8 VSS 0.00452325f
c5 9 VSS 0.00121364f
c6 10 VSS 0.000899441f
c7 11 VSS 0.0065426f
c8 12 VSS 0.00658108f
c9 13 VSS 0.00741325f
c10 14 VSS 0.0021483f
c11 15 VSS 0.00201609f
c12 16 VSS 0.0034704f
c13 17 VSS 0.0034704f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 36 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r6 32 33 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2700 $Y2=0.2160
r7 10 32 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1865 $X2=0.2700 $Y2=0.1980
r8 15 31 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2815 $Y2=0.2340
r9 15 33 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2700 $Y2=0.2160
r10 12 17 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3130 $Y=0.2340 $X2=0.3510 $Y2=0.2340
r11 12 31 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3130
+ $Y=0.2340 $X2=0.2815 $Y2=0.2340
r12 17 30 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.2045
r13 29 30 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1660 $X2=0.3510 $Y2=0.2045
r14 28 29 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1475 $X2=0.3510 $Y2=0.1660
r15 28 27 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1475 $X2=0.3510 $Y2=0.1455
r16 26 27 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1455
r17 25 26 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1060 $X2=0.3510 $Y2=0.1350
r18 13 16 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0655 $X2=0.3510 $Y2=0.0360
r19 13 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0655 $X2=0.3510 $Y2=0.1060
r20 16 24 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0360 $X2=0.3130 $Y2=0.0360
r21 11 14 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2815 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r22 11 24 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2815
+ $Y=0.0360 $X2=0.3130 $Y2=0.0360
r23 9 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0720
r24 9 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0360
r25 1 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0720
r26 21 19 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r27 1 19 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r28 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r29 20 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_OR3x2_ASAP7_75t_R%NET61 VSS 12 13 60 61 63 65 3 17 18 16 4 14 5 15 1
+ 20 19 23 21 24 22
c1 1 VSS 0.00711387f
c2 3 VSS 0.00918298f
c3 4 VSS 0.00714464f
c4 5 VSS 0.009944f
c5 12 VSS 0.0805742f
c6 13 VSS 0.080789f
c7 14 VSS 0.00584915f
c8 15 VSS 0.00665294f
c9 16 VSS 0.00491433f
c10 17 VSS 0.0192549f
c11 18 VSS 0.019861f
c12 19 VSS 0.00241569f
c13 20 VSS 0.00243553f
c14 21 VSS 0.001059f
c15 22 VSS 0.00231486f
c16 23 VSS 0.000174069f
c17 24 VSS 0.00259829f
r1 65 64 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 16 64 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 63 62 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r4 14 62 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r5 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 5 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 15 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 60 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r10 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r11 5 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r12 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 54 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 53 54 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 52 53 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 51 52 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 50 51 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 18 24 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2100 $Y=0.2340 $X2=0.2310 $Y2=0.2340
r19 18 50 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2100
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r20 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r21 46 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r22 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r23 44 45 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r24 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r25 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r26 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r27 40 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r28 17 22 3.24787 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2100 $Y=0.0360 $X2=0.2310 $Y2=0.0360
r29 17 40 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2100
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 24 39 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2310 $Y=0.2340 $X2=0.2310 $Y2=0.2125
r31 22 37 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2310 $Y=0.0360 $X2=0.2310 $Y2=0.0575
r32 38 39 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2310
+ $Y=0.1920 $X2=0.2310 $Y2=0.2125
r33 20 23 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2310 $Y=0.1640 $X2=0.2310 $Y2=0.1350
r34 20 38 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2310
+ $Y=0.1640 $X2=0.2310 $Y2=0.1920
r35 36 37 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2310
+ $Y=0.0780 $X2=0.2310 $Y2=0.0575
r36 19 23 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2310 $Y=0.1060 $X2=0.2310 $Y2=0.1350
r37 19 36 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2310
+ $Y=0.1060 $X2=0.2310 $Y2=0.0780
r38 23 33 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2310 $Y=0.1350 $X2=0.2505 $Y2=0.1350
r39 13 31 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r40 21 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2700 $Y=0.1350
+ $X2=0.2700 $Y2=0.1350
r41 21 33 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2505 $Y2=0.1350
r42 29 31 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r43 28 29 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r44 27 28 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2555 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r45 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r46 1 26 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r47 1 27 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r48 12 26 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r49 12 27 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r50 4 16 1e-05
r51 3 14 1e-05
.ends


*
.SUBCKT OR3x2_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM1@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM12_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM1@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR3x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR3x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR3x2_ASAP7_75t_R%NET67 VSS N_MM11_s N_MM10_d N_NET67_1
+ PM_OR3x2_ASAP7_75t_R%NET67
cc_1 N_NET67_1 N_MM12_g 0.017189f
cc_2 N_NET67_1 N_MM13_g 0.0173141f
x_PM_OR3x2_ASAP7_75t_R%NET66 VSS N_MM10_s N_MM8_d N_NET66_1
+ PM_OR3x2_ASAP7_75t_R%NET66
cc_3 N_NET66_1 N_MM13_g 0.0173501f
cc_4 N_NET66_1 N_MM14_g 0.017378f
x_PM_OR3x2_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR3x2_ASAP7_75t_R%noxref_10
cc_5 N_noxref_10_1 N_MM12_g 0.00162755f
cc_6 N_noxref_10_1 N_NET61_14 0.0381021f
x_PM_OR3x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR3x2_ASAP7_75t_R%noxref_12
cc_7 N_noxref_12_1 N_MM1@2_g 0.00145974f
cc_8 N_noxref_12_1 N_Y_7 0.000830352f
x_PM_OR3x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_OR3x2_ASAP7_75t_R%noxref_13
cc_9 N_noxref_13_1 N_MM1@2_g 0.00146677f
cc_10 N_noxref_13_1 N_Y_8 0.000832578f
cc_11 N_noxref_13_1 N_noxref_12_1 0.00177749f
x_PM_OR3x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR3x2_ASAP7_75t_R%noxref_11
cc_12 N_noxref_11_1 N_MM12_g 0.0016363f
cc_13 N_noxref_11_1 N_NET61_16 0.0380045f
cc_14 N_noxref_11_1 N_noxref_10_1 0.00179378f
x_PM_OR3x2_ASAP7_75t_R%C VSS C N_MM14_g N_C_4 N_C_1 PM_OR3x2_ASAP7_75t_R%C
cc_15 N_MM14_g N_B_1 0.00124419f
cc_16 N_C_4 N_B_4 0.00475331f
cc_17 N_MM14_g N_MM13_g 0.00612829f
x_PM_OR3x2_ASAP7_75t_R%A VSS A N_MM12_g N_A_1 N_A_4 PM_OR3x2_ASAP7_75t_R%A
x_PM_OR3x2_ASAP7_75t_R%B VSS B N_MM13_g N_B_1 N_B_4 PM_OR3x2_ASAP7_75t_R%B
cc_18 N_B_1 N_A_1 0.00119683f
cc_19 N_B_4 N_A_4 0.00483114f
cc_20 N_MM13_g N_MM12_g 0.00626621f
x_PM_OR3x2_ASAP7_75t_R%Y VSS Y N_MM1_d N_MM1@2_d N_MM0_d N_MM0@2_d N_Y_7 N_Y_1
+ N_Y_13 N_Y_15 N_Y_14 N_Y_9 N_Y_2 N_Y_10 N_Y_8 PM_OR3x2_ASAP7_75t_R%Y
cc_21 N_Y_7 N_NET61_20 0.000486851f
cc_22 N_Y_7 N_NET61_19 0.000495053f
cc_23 N_Y_1 N_NET61_1 0.000955038f
cc_24 N_Y_13 N_NET61_21 0.00105593f
cc_25 N_Y_15 N_NET61_24 0.00139478f
cc_26 N_Y_14 N_NET61_22 0.00140944f
cc_27 N_Y_9 N_NET61_21 0.00146505f
cc_28 N_Y_2 N_MM1@2_g 0.0021658f
cc_29 N_Y_1 N_MM1@2_g 0.0021871f
cc_30 N_Y_9 N_NET61_19 0.00398473f
cc_31 N_Y_10 N_NET61_20 0.00402291f
cc_32 N_Y_8 N_NET61_1 0.00444679f
cc_33 N_Y_8 N_MM1@2_g 0.0300788f
cc_34 N_Y_7 N_MM1_g 0.0371838f
cc_35 N_Y_7 N_MM1@2_g 0.0697331f
x_PM_OR3x2_ASAP7_75t_R%NET61 VSS N_MM1_g N_MM1@2_g N_MM13_d N_MM14_d N_MM12_d
+ N_MM11_d N_NET61_3 N_NET61_17 N_NET61_18 N_NET61_16 N_NET61_4 N_NET61_14
+ N_NET61_5 N_NET61_15 N_NET61_1 N_NET61_20 N_NET61_19 N_NET61_23 N_NET61_21
+ N_NET61_24 N_NET61_22 PM_OR3x2_ASAP7_75t_R%NET61
cc_36 N_NET61_3 N_A_1 0.00063074f
cc_37 N_NET61_17 N_A_4 0.0012248f
cc_38 N_NET61_18 N_A_4 0.00139015f
cc_39 N_NET61_3 N_MM12_g 0.00152157f
cc_40 N_NET61_16 N_A_1 0.0016622f
cc_41 N_NET61_4 N_MM12_g 0.00189543f
cc_42 N_NET61_3 N_A_4 0.00428059f
cc_43 N_NET61_16 N_MM12_g 0.0155189f
cc_44 N_NET61_14 N_MM12_g 0.0553769f
cc_45 N_NET61_5 N_MM13_g 0.00151827f
cc_46 N_NET61_15 N_B_1 0.000729046f
cc_47 N_NET61_17 N_B_4 0.00112319f
cc_48 N_NET61_18 N_B_4 0.00140419f
cc_49 N_NET61_5 N_B_4 0.00323778f
cc_50 N_NET61_15 N_MM13_g 0.0360524f
cc_51 N_NET61_1 N_MM14_g 0.000452288f
cc_52 N_NET61_5 N_MM14_g 0.00187366f
cc_53 N_NET61_17 N_MM14_g 0.000909776f
cc_54 N_NET61_18 N_C_4 0.0010973f
cc_55 N_NET61_15 N_C_1 0.00122912f
cc_56 N_MM1_g N_MM14_g 0.00162654f
cc_57 N_NET61_20 N_C_4 0.00174616f
cc_58 N_NET61_19 N_C_4 0.00176748f
cc_59 N_NET61_23 N_C_4 0.00696864f
cc_60 N_NET61_15 N_MM14_g 0.0368551f
*END of OR3x2_ASAP7_75t_R.pxi
.ENDS
** Design:	OR3x4_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR3x4_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR3x4_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR3x4_ASAP7_75t_R%NET66 VSS 2 3 1
c1 1 VSS 0.000959845f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR3x4_ASAP7_75t_R%NET67 VSS 2 3 1
c1 1 VSS 0.000969517f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR3x4_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0422897f
.ends

.subckt PM_OR3x4_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0422896f
.ends

.subckt PM_OR3x4_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00492674f
.ends

.subckt PM_OR3x4_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.00482733f
.ends

.subckt PM_OR3x4_ASAP7_75t_R%C VSS 7 3 4 1
c1 1 VSS 0.00666351f
c2 3 VSS 0.0830636f
c3 4 VSS 0.00457032f
r1 7 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.0980
r2 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 7 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_OR3x4_ASAP7_75t_R%B VSS 6 3 1 4
c1 1 VSS 0.00554724f
c2 3 VSS 0.045934f
c3 4 VSS 0.00402754f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_OR3x4_ASAP7_75t_R%A VSS 6 3 1 4
c1 1 VSS 0.00268139f
c2 3 VSS 0.0429861f
c3 4 VSS 0.0122266f
r1 6 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r2 3 1 7.10798 $w=1.13765e-07 $l=5e-10 $layer=LIG $thickness=5.17209e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1355
r3 6 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1355
.ends

.subckt PM_OR3x4_ASAP7_75t_R%Y VSS 48 34 35 43 44 58 59 62 63 13 1 2 14 15 16
+ 27 17 26 4 3 18
c1 1 VSS 0.00833009f
c2 2 VSS 0.00829139f
c3 3 VSS 0.00850561f
c4 4 VSS 0.00848692f
c5 13 VSS 0.00453008f
c6 14 VSS 0.00442704f
c7 15 VSS 0.00450753f
c8 16 VSS 0.00441415f
c9 17 VSS 0.00125987f
c10 18 VSS 0.00089423f
c11 19 VSS 0.00912901f
c12 20 VSS 0.00910543f
c13 21 VSS 0.0010654f
c14 22 VSS 0.0010654f
c15 23 VSS 0.00641946f
c16 24 VSS 0.00641946f
c17 25 VSS 0.00721591f
c18 26 VSS 0.0023082f
c19 27 VSS 0.00209357f
c20 28 VSS 0.00249529f
c21 29 VSS 0.00249529f
c22 30 VSS 0.00344782f
c23 31 VSS 0.00344782f
r1 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 62 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 54 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.1980
r6 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r7 4 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r8 16 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r9 58 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r10 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2700 $Y2=0.2160
r11 18 54 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1865 $X2=0.2700 $Y2=0.1980
r12 4 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.1980
r13 27 51 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2815 $Y2=0.2340
r14 27 55 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.2700 $Y2=0.2160
r15 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1980 $X2=0.3780 $Y2=0.2160
r16 22 52 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.1865 $X2=0.3780 $Y2=0.1980
r17 20 29 10.829 $w=1.38738e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3265 $Y=0.2340 $X2=0.3780 $Y2=0.2340
r18 20 51 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3265
+ $Y=0.2340 $X2=0.2815 $Y2=0.2340
r19 29 53 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3780 $Y2=0.2160
r20 24 31 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4185 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r21 24 29 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4185 $Y=0.2340 $X2=0.3780 $Y2=0.2340
r22 31 50 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4590 $Y2=0.2045
r23 49 50 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1660 $X2=0.4590 $Y2=0.2045
r24 48 49 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1660
r25 48 47 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1455
r26 46 47 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1455
r27 45 46 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1060 $X2=0.4590 $Y2=0.1350
r28 25 30 5.22999 $w=1.59898e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0655 $X2=0.4590 $Y2=0.0360
r29 25 45 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0655 $X2=0.4590 $Y2=0.1060
r30 44 42 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r31 3 42 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r32 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r33 43 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r34 3 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0720
r35 23 28 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4185 $Y=0.0360 $X2=0.3780 $Y2=0.0360
r36 23 30 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4185 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r37 21 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0540 $X2=0.3780 $Y2=0.0720
r38 21 28 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0540 $X2=0.3780 $Y2=0.0360
r39 28 38 10.829 $w=1.38738e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3780 $Y=0.0360 $X2=0.3265 $Y2=0.0360
r40 19 26 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2815 $Y=0.0360 $X2=0.2700 $Y2=0.0360
r41 19 38 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2815
+ $Y=0.0360 $X2=0.3265 $Y2=0.0360
r42 17 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0720
r43 17 26 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0360
r44 1 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0720
r45 35 33 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r46 1 33 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r47 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r48 34 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_OR3x4_ASAP7_75t_R%NET61 VSS 12 13 14 15 78 79 81 83 18 3 19 20 4 16
+ 5 17 1 21 22 25 26 24 23
c1 1 VSS 0.0160557f
c2 3 VSS 0.01029f
c3 4 VSS 0.0082878f
c4 5 VSS 0.00991204f
c5 12 VSS 0.0806261f
c6 13 VSS 0.080358f
c7 14 VSS 0.080089f
c8 15 VSS 0.0806623f
c9 16 VSS 0.0088522f
c10 17 VSS 0.00938076f
c11 18 VSS 0.00790631f
c12 19 VSS 0.0218407f
c13 20 VSS 0.0224082f
c14 21 VSS 0.00294609f
c15 22 VSS 0.00299394f
c16 23 VSS 0.00141518f
c17 24 VSS 0.0028126f
c18 25 VSS 0.000252496f
c19 26 VSS 0.00250631f
r1 83 82 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 18 82 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 81 80 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r4 16 80 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r5 79 77 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r6 5 77 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r7 17 5 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r8 78 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r9 4 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r10 3 66 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r11 5 60 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r12 74 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r13 72 75 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r14 71 72 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.0810 $Y2=0.2340
r15 70 71 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r16 69 70 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r17 68 69 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.2340 $X2=0.1620 $Y2=0.2340
r18 20 26 3.36447 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2105 $Y=0.2340 $X2=0.2320 $Y2=0.2340
r19 20 68 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2105
+ $Y=0.2340 $X2=0.1890 $Y2=0.2340
r20 66 67 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r21 64 67 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r22 63 64 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r23 62 63 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r24 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r25 59 60 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r26 59 62 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r27 58 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r28 19 24 3.36447 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2105 $Y=0.0360 $X2=0.2320 $Y2=0.0360
r29 19 58 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2105
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r30 26 57 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.2340 $X2=0.2320 $Y2=0.2125
r31 24 55 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.0360 $X2=0.2320 $Y2=0.0575
r32 56 57 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1920 $X2=0.2320 $Y2=0.2125
r33 22 25 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.1640 $X2=0.2320 $Y2=0.1350
r34 22 56 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1640 $X2=0.2320 $Y2=0.1920
r35 54 55 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.0780 $X2=0.2320 $Y2=0.0575
r36 21 25 5.5822 $w=1.45517e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.1060 $X2=0.2320 $Y2=0.1350
r37 21 54 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.1060 $X2=0.2320 $Y2=0.0780
r38 25 49 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2320 $Y=0.1350 $X2=0.2510 $Y2=0.1350
r39 15 47 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r40 14 41 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r41 13 35 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r42 23 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2700 $Y=0.1350
+ $X2=0.2700 $Y2=0.1350
r43 23 49 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2510 $Y2=0.1350
r44 45 47 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r45 44 45 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r46 42 44 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r47 41 42 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r48 39 41 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r49 38 39 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r50 36 38 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r51 35 36 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r52 33 35 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r53 32 33 2.36289 $w=1.53e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.2805
+ $Y=0.1350 $X2=0.2845 $Y2=0.1350
r54 31 32 6.20259 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2700 $Y=0.1350 $X2=0.2805 $Y2=0.1350
r55 30 31 6.20259 $w=1.53e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2595 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r56 29 30 2.36289 $w=1.53e-08 $l=4e-09 $layer=LIG $thickness=4.8e-08 $X=0.2555
+ $Y=0.1350 $X2=0.2595 $Y2=0.1350
r57 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r58 1 28 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r59 1 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r60 12 28 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2325 $Y2=0.1350
r61 12 29 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2555 $Y2=0.1350
r62 4 18 1e-05
r63 3 16 1e-05
.ends


*
.SUBCKT OR3x4_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM12 N_MM12_d N_MM12_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM13_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@4 N_MM1@4_d N_MM0@4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@3 N_MM1@3_d N_MM0@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 N_MM1@2_d N_MM0@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM12_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM13_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@4 N_MM0@4_d N_MM0@4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@3 N_MM0@3_d N_MM0@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0@2 N_MM0@2_d N_MM0@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR3x4_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR3x4_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR3x4_ASAP7_75t_R%NET66 VSS N_MM10_s N_MM8_d N_NET66_1
+ PM_OR3x4_ASAP7_75t_R%NET66
cc_1 N_NET66_1 N_MM13_g 0.0173496f
cc_2 N_NET66_1 N_MM14_g 0.017379f
x_PM_OR3x4_ASAP7_75t_R%NET67 VSS N_MM11_s N_MM10_d N_NET67_1
+ PM_OR3x4_ASAP7_75t_R%NET67
cc_3 N_NET67_1 N_MM12_g 0.0171923f
cc_4 N_NET67_1 N_MM13_g 0.0173186f
x_PM_OR3x4_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_OR3x4_ASAP7_75t_R%noxref_13
cc_5 N_noxref_13_1 N_MM0@2_g 0.00145985f
cc_6 N_noxref_13_1 N_Y_16 0.000830636f
cc_7 N_noxref_13_1 N_noxref_12_1 0.00178875f
x_PM_OR3x4_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR3x4_ASAP7_75t_R%noxref_12
cc_8 N_noxref_12_1 N_MM0@2_g 0.00145591f
cc_9 N_noxref_12_1 N_Y_14 0.00083008f
x_PM_OR3x4_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_OR3x4_ASAP7_75t_R%noxref_11
cc_10 N_noxref_11_1 N_MM12_g 0.00163597f
cc_11 N_noxref_11_1 N_NET61_4 0.000542124f
cc_12 N_noxref_11_1 N_NET61_18 0.0374655f
cc_13 N_noxref_11_1 N_noxref_10_1 0.00179311f
x_PM_OR3x4_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_OR3x4_ASAP7_75t_R%noxref_10
cc_14 N_noxref_10_1 N_MM12_g 0.00162921f
cc_15 N_noxref_10_1 N_NET61_3 0.000538521f
cc_16 N_noxref_10_1 N_NET61_16 0.0375705f
x_PM_OR3x4_ASAP7_75t_R%C VSS C N_MM14_g N_C_4 N_C_1 PM_OR3x4_ASAP7_75t_R%C
cc_17 N_MM14_g N_B_1 0.00126993f
cc_18 N_C_4 N_B_4 0.0047579f
cc_19 N_MM14_g N_MM13_g 0.0061471f
x_PM_OR3x4_ASAP7_75t_R%B VSS B N_MM13_g N_B_1 N_B_4 PM_OR3x4_ASAP7_75t_R%B
cc_20 N_B_1 N_A_1 0.00127096f
cc_21 N_B_4 N_A_4 0.00482282f
cc_22 N_MM13_g N_MM12_g 0.00626622f
x_PM_OR3x4_ASAP7_75t_R%A VSS A N_MM12_g N_A_1 N_A_4 PM_OR3x4_ASAP7_75t_R%A
x_PM_OR3x4_ASAP7_75t_R%Y VSS Y N_MM1_d N_MM1@4_d N_MM1@3_d N_MM1@2_d N_MM0@3_d
+ N_MM0@2_d N_MM0_d N_MM0@4_d N_Y_13 N_Y_1 N_Y_2 N_Y_14 N_Y_15 N_Y_16 N_Y_27
+ N_Y_17 N_Y_26 N_Y_4 N_Y_3 N_Y_18 PM_OR3x4_ASAP7_75t_R%Y
cc_23 N_Y_13 N_NET61_1 0.00121685f
cc_24 N_Y_13 N_NET61_26 0.000295081f
cc_25 N_Y_13 N_NET61_24 0.000311812f
cc_26 N_Y_1 N_NET61_21 0.000519154f
cc_27 N_Y_2 N_NET61_22 0.000608725f
cc_28 N_Y_14 N_MM0@2_g 0.0675306f
cc_29 N_Y_15 N_MM0@4_g 0.0307341f
cc_30 N_Y_16 N_MM0@2_g 0.0307463f
cc_31 N_Y_1 N_NET61_1 0.000895121f
cc_32 N_Y_27 N_NET61_26 0.0012395f
cc_33 N_Y_17 N_NET61_23 0.00128363f
cc_34 N_Y_26 N_NET61_24 0.00149893f
cc_35 N_Y_4 N_MM0@2_g 0.00174849f
cc_36 N_Y_3 N_MM0@2_g 0.00176354f
cc_37 N_Y_2 N_MM0@4_g 0.00221205f
cc_38 N_Y_1 N_MM0@4_g 0.00221819f
cc_39 N_Y_18 N_NET61_22 0.00391206f
cc_40 N_Y_17 N_NET61_21 0.00399448f
cc_41 N_Y_16 N_NET61_1 0.00941276f
cc_42 N_Y_13 N_MM0_g 0.0368446f
cc_43 N_Y_14 N_MM0@3_g 0.0368909f
cc_44 N_Y_13 N_MM0@4_g 0.0685322f
x_PM_OR3x4_ASAP7_75t_R%NET61 VSS N_MM0_g N_MM0@4_g N_MM0@3_g N_MM0@2_g N_MM13_d
+ N_MM14_d N_MM12_d N_MM11_d N_NET61_18 N_NET61_3 N_NET61_19 N_NET61_20
+ N_NET61_4 N_NET61_16 N_NET61_5 N_NET61_17 N_NET61_1 N_NET61_21 N_NET61_22
+ N_NET61_25 N_NET61_26 N_NET61_24 N_NET61_23 PM_OR3x4_ASAP7_75t_R%NET61
cc_45 N_NET61_18 N_MM12_g 0.0159818f
cc_46 N_NET61_3 N_A_1 0.00063074f
cc_47 N_NET61_19 N_A_4 0.00129408f
cc_48 N_NET61_20 N_A_4 0.0013841f
cc_49 N_NET61_3 N_MM12_g 0.00152157f
cc_50 N_NET61_18 N_A_1 0.0016622f
cc_51 N_NET61_4 N_MM12_g 0.00190233f
cc_52 N_NET61_3 N_A_4 0.00429695f
cc_53 N_NET61_16 N_MM12_g 0.0549108f
cc_54 N_NET61_4 N_MM13_g 0.000288101f
cc_55 N_NET61_5 N_MM13_g 0.0015181f
cc_56 N_NET61_17 N_B_1 0.000862656f
cc_57 N_NET61_19 N_B_4 0.00122963f
cc_58 N_NET61_20 N_B_4 0.00140586f
cc_59 N_NET61_5 N_B_4 0.00325291f
cc_60 N_NET61_17 N_MM13_g 0.035808f
cc_61 N_NET61_1 N_MM14_g 0.0004329f
cc_62 N_NET61_5 N_MM14_g 0.00185253f
cc_63 N_NET61_19 N_MM14_g 0.00100552f
cc_64 N_NET61_20 N_C_4 0.00115907f
cc_65 N_NET61_17 N_C_1 0.00120594f
cc_66 N_MM0_g N_MM14_g 0.00164922f
cc_67 N_NET61_21 N_C_4 0.00171999f
cc_68 N_NET61_22 N_C_4 0.00178732f
cc_69 N_NET61_25 N_C_4 0.00711731f
cc_70 N_NET61_17 N_MM14_g 0.0368393f
*END of OR3x4_ASAP7_75t_R.pxi
.ENDS
** Design:	OR4x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR4x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR4x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR4x1_ASAP7_75t_R%PD2 VSS 2 3 1
c1 1 VSS 0.000901995f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_OR4x1_ASAP7_75t_R%PD1 VSS 2 3 1
c1 1 VSS 0.00092577f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_OR4x1_ASAP7_75t_R%PD3 VSS 2 3 1
c1 1 VSS 0.000920454f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR4x1_ASAP7_75t_R%Y VSS 13 24 7 2 8 1 10 9
c1 1 VSS 0.00814826f
c2 2 VSS 0.00943056f
c3 7 VSS 0.00384042f
c4 8 VSS 0.00380006f
c5 9 VSS 0.0040483f
c6 10 VSS 0.0051568f
c7 11 VSS 0.00640713f
r1 24 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 8 23 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 20 21 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 11 19 9.42983 $w=1.3989e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.1885
r6 11 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 18 19 16.4399 $w=1.3e-08 $l=7.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1180 $X2=0.0270 $Y2=0.1885
r8 17 18 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0750 $X2=0.0270 $Y2=0.1180
r9 9 16 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0555 $X2=0.0270 $Y2=0.0360
r10 9 17 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0555 $X2=0.0270 $Y2=0.0750
r11 10 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r12 10 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0405 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r13 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r14 13 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r15 7 12 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r16 2 8 1e-05
r17 1 7 1e-05
.ends

.subckt PM_OR4x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0419663f
.ends

.subckt PM_OR4x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00529001f
.ends

.subckt PM_OR4x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00474848f
.ends

.subckt PM_OR4x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00466055f
.ends

.subckt PM_OR4x1_ASAP7_75t_R%D VSS 8 3 1 4
c1 1 VSS 0.00658504f
c2 3 VSS 0.0835872f
c3 4 VSS 0.00925971f
r1 8 4 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1160
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
.ends

.subckt PM_OR4x1_ASAP7_75t_R%A VSS 8 3 4 1
c1 1 VSS 0.00674108f
c2 3 VSS 0.045663f
c3 4 VSS 0.0049526f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_OR4x1_ASAP7_75t_R%C VSS 10 3 1 4
c1 1 VSS 0.00587081f
c2 3 VSS 0.0464154f
c3 4 VSS 0.00761069f
r1 10 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1160
r2 4 9 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0950 $X2=0.1890 $Y2=0.1160
r3 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_OR4x1_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00527185f
c2 3 VSS 0.0458297f
c3 4 VSS 0.00733598f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_OR4x1_ASAP7_75t_R%NET12 VSS 12 47 48 51 52 60 1 20 3 13 16 18 4 5 14
+ 22 15 19 21
c1 1 VSS 0.00321192f
c2 3 VSS 0.00998924f
c3 4 VSS 0.00995948f
c4 5 VSS 0.00631962f
c5 12 VSS 0.0800411f
c6 13 VSS 0.00493927f
c7 14 VSS 0.00492117f
c8 15 VSS 0.00323355f
c9 16 VSS 0.00129131f
c10 17 VSS 0.000792523f
c11 18 VSS 0.0212618f
c12 19 VSS 0.00541257f
c13 20 VSS 0.00133637f
c14 21 VSS 0.0026718f
c15 22 VSS 0.00636852f
c16 23 VSS 0.00343605f
r1 15 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 60 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 5 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r4 57 58 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.2340 $X2=0.3375 $Y2=0.2340
r5 22 55 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3510 $Y2=0.2125
r6 22 58 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.2340 $X2=0.3375 $Y2=0.2340
r7 54 55 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.2125
r8 53 54 15.6237 $w=1.3e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0680 $X2=0.3510 $Y2=0.1350
r9 19 23 2.89809 $w=1.75231e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0555 $X2=0.3510 $Y2=0.0360
r10 19 53 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0555 $X2=0.3510 $Y2=0.0680
r11 52 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r12 4 50 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r13 14 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r14 51 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r15 48 46 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r16 3 46 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0675 $X2=0.1765 $Y2=0.0675
r17 13 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r18 47 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r19 23 44 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3260 $Y2=0.0360
r20 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r21 3 34 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0675
+ $X2=0.1620 $Y2=0.0360
r22 43 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3080
+ $Y=0.0360 $X2=0.3260 $Y2=0.0360
r23 42 43 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3080 $Y2=0.0360
r24 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r25 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r26 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r27 38 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2565 $Y2=0.0360
r28 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r29 36 37 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r30 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r31 34 35 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r32 33 34 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r33 32 33 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1485 $Y2=0.0360
r34 18 21 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1215 $Y=0.0360 $X2=0.1080 $Y2=0.0360
r35 18 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r36 17 31 3.36689 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0555 $X2=0.1080 $Y2=0.0750
r37 17 21 2.89809 $w=1.75231e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0555 $X2=0.1080 $Y2=0.0360
r38 30 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0750 $X2=0.1080 $Y2=0.0750
r39 20 29 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0750 $X2=0.0810 $Y2=0.0950
r40 20 30 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0750 $X2=0.0945 $Y2=0.0750
r41 16 27 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1350
r42 16 29 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.0950
r43 12 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r44 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends


*
.SUBCKT OR4x1_ASAP7_75t_R VSS VDD D C B A
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
*
*

MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM1_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM0_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR4x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR4x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR4x1_ASAP7_75t_R%PD2 VSS N_MM5_d N_MM6_s N_PD2_1 PM_OR4x1_ASAP7_75t_R%PD2
cc_1 N_PD2_1 N_MM2_g 0.017332f
cc_2 N_PD2_1 N_MM1_g 0.0173902f
x_PM_OR4x1_ASAP7_75t_R%PD1 VSS N_MM6_d N_MM7_s N_PD1_1 PM_OR4x1_ASAP7_75t_R%PD1
cc_3 N_PD1_1 N_MM1_g 0.0172205f
cc_4 N_PD1_1 N_MM0_g 0.0172362f
x_PM_OR4x1_ASAP7_75t_R%PD3 VSS N_MM4_d N_MM5_s N_PD3_1 PM_OR4x1_ASAP7_75t_R%PD3
cc_5 N_PD3_1 N_MM3_g 0.0171868f
cc_6 N_PD3_1 N_MM2_g 0.0172968f
x_PM_OR4x1_ASAP7_75t_R%Y VSS N_MM9_d N_MM8_d N_Y_7 N_Y_2 N_Y_8 N_Y_1 N_Y_10
+ N_Y_9 PM_OR4x1_ASAP7_75t_R%Y
cc_7 N_Y_7 N_NET12_21 0.000402768f
cc_8 N_Y_7 N_NET12_1 0.000943755f
cc_9 N_Y_2 N_MM9_g 0.00101715f
cc_10 N_Y_8 N_NET12_1 0.00132636f
cc_11 N_Y_1 N_MM9_g 0.00140727f
cc_12 N_Y_10 N_NET12_20 0.00202682f
cc_13 N_Y_9 N_NET12_16 0.00450827f
cc_14 N_Y_8 N_MM9_g 0.0153936f
cc_15 N_Y_7 N_MM9_g 0.0550797f
x_PM_OR4x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_OR4x1_ASAP7_75t_R%noxref_14
cc_16 N_noxref_14_1 N_NET12_14 0.00131439f
cc_17 N_noxref_14_1 N_MM0_g 0.00145635f
x_PM_OR4x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_OR4x1_ASAP7_75t_R%noxref_15
cc_18 N_noxref_15_1 N_NET12_15 0.0379125f
cc_19 N_noxref_15_1 N_MM0_g 0.00145893f
cc_20 N_noxref_15_1 N_noxref_14_1 0.00178178f
x_PM_OR4x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR4x1_ASAP7_75t_R%noxref_12
cc_21 N_noxref_12_1 N_MM9_g 0.00146012f
cc_22 N_noxref_12_1 N_Y_7 0.0384656f
x_PM_OR4x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_OR4x1_ASAP7_75t_R%noxref_13
cc_23 N_noxref_13_1 N_MM9_g 0.00144324f
cc_24 N_noxref_13_1 N_Y_8 0.0385403f
cc_25 N_noxref_13_1 N_noxref_12_1 0.00177728f
x_PM_OR4x1_ASAP7_75t_R%D VSS D N_MM3_g N_D_1 N_D_4 PM_OR4x1_ASAP7_75t_R%D
cc_26 N_MM3_g N_NET12_1 0.000478676f
cc_27 N_MM3_g N_NET12_20 0.000491561f
cc_28 N_MM3_g N_NET12_3 0.00160471f
cc_29 N_D_1 N_NET12_13 0.000947031f
cc_30 N_MM3_g N_MM9_g 0.00165839f
cc_31 N_D_4 N_NET12_16 0.00339956f
cc_32 N_MM3_g N_NET12_13 0.0369472f
x_PM_OR4x1_ASAP7_75t_R%A VSS A N_MM0_g N_A_4 N_A_1 PM_OR4x1_ASAP7_75t_R%A
cc_33 N_A_4 N_NET12_22 0.000512604f
cc_34 N_A_1 N_NET12_5 0.00095371f
cc_35 N_A_4 N_NET12_18 0.00111326f
cc_36 N_MM0_g N_NET12_4 0.00115268f
cc_37 N_A_1 N_NET12_15 0.00140465f
cc_38 N_MM0_g N_NET12_5 0.00168175f
cc_39 N_MM0_g N_NET12_15 0.0154213f
cc_40 N_A_4 N_NET12_19 0.00823828f
cc_41 N_MM0_g N_NET12_14 0.0549872f
cc_42 N_A_1 N_B_1 0.00111017f
cc_43 N_MM0_g N_MM1_g 0.00520266f
cc_44 N_A_4 N_B_4 0.00652428f
x_PM_OR4x1_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 N_C_4 PM_OR4x1_ASAP7_75t_R%C
cc_45 N_C_1 N_NET12_13 0.000686456f
cc_46 N_MM2_g N_NET12_3 0.00122337f
cc_47 N_C_4 N_NET12_18 0.00126152f
cc_48 N_C_4 N_NET12_3 0.00213439f
cc_49 N_MM2_g N_NET12_13 0.0356871f
cc_50 N_C_1 N_D_4 0.00109338f
cc_51 N_MM2_g N_MM3_g 0.00522176f
cc_52 N_C_4 N_D_4 0.00648274f
x_PM_OR4x1_ASAP7_75t_R%B VSS B N_MM1_g N_B_1 N_B_4 PM_OR4x1_ASAP7_75t_R%B
cc_53 N_MM1_g N_NET12_4 0.0015069f
cc_54 N_MM1_g N_NET12_5 0.000348923f
cc_55 N_B_1 N_NET12_14 0.000635276f
cc_56 N_B_4 N_NET12_18 0.00119185f
cc_57 N_B_4 N_NET12_4 0.00232552f
cc_58 N_MM1_g N_NET12_14 0.0358341f
cc_59 N_B_1 N_C_1 0.00113301f
cc_60 N_MM1_g N_MM2_g 0.00543468f
cc_61 N_B_4 N_C_4 0.00752106f
x_PM_OR4x1_ASAP7_75t_R%NET12 VSS N_MM9_g N_MM3_d N_MM2_d N_MM1_d N_MM0_d
+ N_MM7_d N_NET12_1 N_NET12_20 N_NET12_3 N_NET12_13 N_NET12_16 N_NET12_18
+ N_NET12_4 N_NET12_5 N_NET12_14 N_NET12_22 N_NET12_15 N_NET12_19 N_NET12_21
+ PM_OR4x1_ASAP7_75t_R%NET12
*END of OR4x1_ASAP7_75t_R.pxi
.ENDS
** Design:	OR4x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR4x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR4x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR4x2_ASAP7_75t_R%PD2 VSS 2 3 1
c1 1 VSS 0.000885038f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_OR4x2_ASAP7_75t_R%PD3 VSS 2 3 1
c1 1 VSS 0.000937936f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_OR4x2_ASAP7_75t_R%PD1 VSS 2 3 1
c1 1 VSS 0.000926497f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3240 $Y2=0.2025
.ends

.subckt PM_OR4x2_ASAP7_75t_R%D VSS 8 3 4 1
c1 1 VSS 0.00696838f
c2 3 VSS 0.0836575f
c3 4 VSS 0.009548f
r1 8 4 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1160
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
.ends

.subckt PM_OR4x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.042342f
.ends

.subckt PM_OR4x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0423423f
.ends

.subckt PM_OR4x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0419692f
.ends

.subckt PM_OR4x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00524455f
.ends

.subckt PM_OR4x2_ASAP7_75t_R%A VSS 8 3 4 1
c1 1 VSS 0.00679103f
c2 3 VSS 0.0455839f
c3 4 VSS 0.00491992f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.0980
r2 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
.ends

.subckt PM_OR4x2_ASAP7_75t_R%Y VSS 21 16 17 28 29 7 10 9 1 2 8
c1 1 VSS 0.0101275f
c2 2 VSS 0.0118825f
c3 7 VSS 0.00460027f
c4 8 VSS 0.00455314f
c5 9 VSS 0.00743521f
c6 10 VSS 0.00890164f
c7 11 VSS 0.00970096f
c8 12 VSS 0.00346335f
c9 13 VSS 0.00341205f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r6 11 13 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.2340 $X2=0.0270 $Y2=0.2340
r7 11 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r8 13 23 9.31081 $w=1.48766e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.1870
r9 22 23 10.785 $w=1.3e-08 $l=4.63e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1407 $X2=0.0270 $Y2=0.1870
r10 21 22 2.04041 $w=1.3e-08 $l=8.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1320 $X2=0.0270 $Y2=0.1407
r11 21 20 8.10334 $w=1.3e-08 $l=3.48e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1320 $X2=0.0270 $Y2=0.0972
r12 9 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r13 9 20 10.0855 $w=1.3e-08 $l=4.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0972
r14 10 18 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r15 10 12 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0675 $Y=0.0360 $X2=0.0270 $Y2=0.0360
r16 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r17 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r18 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r20 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_OR4x2_ASAP7_75t_R%C VSS 10 3 1 4
c1 1 VSS 0.00549226f
c2 3 VSS 0.0463396f
c3 4 VSS 0.00788974f
r1 10 9 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1160
r2 4 9 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0935 $X2=0.2430 $Y2=0.1160
r3 3 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_OR4x2_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00564822f
c2 3 VSS 0.0459452f
c3 4 VSS 0.00747878f
r1 8 4 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.0980
r2 3 1 3.49039 $w=1.235e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_OR4x2_ASAP7_75t_R%NET12 VSS 12 13 56 57 60 61 68 20 24 1 3 17 14 21
+ 4 5 15 16 25 23 22 18
c1 1 VSS 0.0067408f
c2 3 VSS 0.00986833f
c3 4 VSS 0.00997315f
c4 5 VSS 0.00651714f
c5 12 VSS 0.0811668f
c6 13 VSS 0.0808638f
c7 14 VSS 0.00639793f
c8 15 VSS 0.00640843f
c9 16 VSS 0.00479342f
c10 17 VSS 0.00210634f
c11 18 VSS 0.00116641f
c12 19 VSS 0.000692014f
c13 20 VSS 0.022596f
c14 21 VSS 0.00873938f
c15 22 VSS 0.000462463f
c16 23 VSS 0.00276576f
c17 24 VSS 0.000904555f
c18 25 VSS 0.00718f
c19 26 VSS 0.00392265f
r1 16 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 68 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 5 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r4 65 66 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r5 25 63 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.4050 $Y2=0.2125
r6 25 66 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.3915 $Y2=0.2340
r7 62 63 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.2125
r8 21 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0575 $X2=0.4050 $Y2=0.0360
r9 21 62 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0575 $X2=0.4050 $Y2=0.1350
r10 61 59 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r11 4 59 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3240 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r12 15 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r13 60 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r14 57 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r15 3 55 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r16 14 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r17 56 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r18 26 53 4.18063 $w=1.48e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.3800 $Y2=0.0360
r19 4 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r20 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r21 52 53 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.0360 $X2=0.3800 $Y2=0.0360
r22 51 52 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0360 $X2=0.3620 $Y2=0.0360
r23 50 51 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3375
+ $Y=0.0360 $X2=0.3510 $Y2=0.0360
r24 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0360 $X2=0.3375 $Y2=0.0360
r25 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3105
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r26 47 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0360 $X2=0.3105 $Y2=0.0360
r27 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2970 $Y2=0.0360
r28 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r29 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2295
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r30 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.2295 $Y2=0.0360
r31 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r32 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r33 20 23 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1755 $Y=0.0360 $X2=0.1620 $Y2=0.0360
r34 20 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1755
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r35 19 24 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0540 $X2=0.1620 $Y2=0.0665
r36 19 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0540 $X2=0.1620 $Y2=0.0360
r37 24 39 3.9716 $w=1.39211e-08 $l=2.51098e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1620 $Y=0.0665 $X2=0.1375 $Y2=0.0720
r38 18 22 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1195 $Y=0.0720 $X2=0.1080 $Y2=0.0720
r39 18 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1195
+ $Y=0.0720 $X2=0.1375 $Y2=0.0720
r40 22 37 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1080 $Y=0.0720 $X2=0.1080 $Y2=0.0935
r41 13 33 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r42 17 35 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1160 $X2=0.1080 $Y2=0.1350
r43 17 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.1160 $X2=0.1080 $Y2=0.0935
r44 31 33 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r45 30 31 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r46 30 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1080 $Y=0.1350
+ $X2=0.1080 $Y2=0.1350
r47 29 30 22.4112 $w=1.13e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r48 12 1 4.17987 $w=1.225e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r49 1 28 4.63801 $w=1.7681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r50 1 29 7.72921 $w=1.666e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r51 12 28 1.08747 $w=2.16729e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r52 12 29 4.17867 $w=1.8386e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT OR4x2_ASAP7_75t_R VSS VDD D C B A Y
*
* VSS VSS
* VDD VDD
* D D
* C C
* B B
* A A
* Y Y
*
*

MM9 N_MM9_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM9@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8@2 N_MM8@2_d N_MM9@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM2_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g N_MM7_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR4x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR4x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR4x2_ASAP7_75t_R%PD2 VSS N_MM6_s N_MM5_d N_PD2_1 PM_OR4x2_ASAP7_75t_R%PD2
cc_1 N_PD2_1 N_MM2_g 0.0173944f
cc_2 N_PD2_1 N_MM6_g 0.0173462f
x_PM_OR4x2_ASAP7_75t_R%PD3 VSS N_MM4_d N_MM5_s N_PD3_1 PM_OR4x2_ASAP7_75t_R%PD3
cc_3 N_PD3_1 N_MM3_g 0.0172359f
cc_4 N_PD3_1 N_MM2_g 0.0172305f
x_PM_OR4x2_ASAP7_75t_R%PD1 VSS N_MM6_d N_MM7_s N_PD1_1 PM_OR4x2_ASAP7_75t_R%PD1
cc_5 N_PD1_1 N_MM6_g 0.0172941f
cc_6 N_PD1_1 N_MM7_g 0.0171621f
x_PM_OR4x2_ASAP7_75t_R%D VSS D N_MM3_g N_D_4 N_D_1 PM_OR4x2_ASAP7_75t_R%D
cc_7 N_MM3_g N_NET12_20 0.000217947f
cc_8 N_MM3_g N_NET12_24 0.000445898f
cc_9 N_MM3_g N_NET12_1 0.000501746f
cc_10 N_MM3_g N_NET12_3 0.001518f
cc_11 N_D_4 N_NET12_17 0.000555002f
cc_12 N_D_1 N_NET12_14 0.00101098f
cc_13 N_MM3_g N_MM9@2_g 0.00165664f
cc_14 N_D_4 N_NET12_1 0.0017007f
cc_15 N_MM3_g N_NET12_14 0.0369389f
x_PM_OR4x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_OR4x2_ASAP7_75t_R%noxref_13
cc_16 N_noxref_13_1 N_MM9_g 0.00146962f
cc_17 N_noxref_13_1 N_Y_8 0.000832311f
cc_18 N_noxref_13_1 N_noxref_12_1 0.00177715f
x_PM_OR4x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_OR4x2_ASAP7_75t_R%noxref_12
cc_19 N_noxref_12_1 N_MM9_g 0.00147219f
cc_20 N_noxref_12_1 N_Y_7 0.000836093f
x_PM_OR4x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_OR4x2_ASAP7_75t_R%noxref_14
cc_21 N_noxref_14_1 N_NET12_15 0.00131488f
cc_22 N_noxref_14_1 N_MM7_g 0.00145726f
x_PM_OR4x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_OR4x2_ASAP7_75t_R%noxref_15
cc_23 N_noxref_15_1 N_NET12_5 0.000506524f
cc_24 N_noxref_15_1 N_NET12_16 0.0374617f
cc_25 N_noxref_15_1 N_MM7_g 0.00145668f
cc_26 N_noxref_15_1 N_noxref_14_1 0.00177642f
x_PM_OR4x2_ASAP7_75t_R%A VSS A N_MM7_g N_A_4 N_A_1 PM_OR4x2_ASAP7_75t_R%A
cc_27 N_MM7_g N_NET12_16 0.0159036f
cc_28 N_A_4 N_NET12_25 0.000572309f
cc_29 N_A_1 N_NET12_5 0.000903332f
cc_30 N_A_4 N_NET12_20 0.0011516f
cc_31 N_MM7_g N_NET12_4 0.00121131f
cc_32 N_A_1 N_NET12_16 0.00145529f
cc_33 N_MM7_g N_NET12_5 0.00167152f
cc_34 N_A_4 N_NET12_21 0.00805736f
cc_35 N_MM7_g N_NET12_15 0.0544921f
cc_36 N_A_1 N_B_1 0.00118768f
cc_37 N_MM7_g N_MM6_g 0.00520938f
cc_38 N_A_4 N_B_4 0.00640562f
x_PM_OR4x2_ASAP7_75t_R%Y VSS Y N_MM9_d N_MM9@2_d N_MM8_d N_MM8@2_d N_Y_7 N_Y_10
+ N_Y_9 N_Y_1 N_Y_2 N_Y_8 PM_OR4x2_ASAP7_75t_R%Y
cc_39 N_Y_7 N_NET12_17 0.00031979f
cc_40 N_Y_7 N_NET12_23 0.000344665f
cc_41 N_Y_7 N_NET12_22 0.000472038f
cc_42 N_Y_7 N_NET12_1 0.000796772f
cc_43 N_Y_10 N_NET12_18 0.000959239f
cc_44 N_Y_9 N_NET12_1 0.00141381f
cc_45 N_Y_1 N_NET12_17 0.00180055f
cc_46 N_Y_2 N_MM9_g 0.00189279f
cc_47 N_Y_1 N_MM9_g 0.00248548f
cc_48 N_Y_10 N_NET12_22 0.00327955f
cc_49 N_Y_8 N_NET12_1 0.00386068f
cc_50 N_Y_8 N_MM9_g 0.0298371f
cc_51 N_Y_7 N_MM9@2_g 0.0371823f
cc_52 N_Y_7 N_MM9_g 0.0693968f
x_PM_OR4x2_ASAP7_75t_R%C VSS C N_MM2_g N_C_1 N_C_4 PM_OR4x2_ASAP7_75t_R%C
cc_53 N_MM2_g N_NET12_3 0.00149016f
cc_54 N_C_1 N_NET12_14 0.000551316f
cc_55 N_C_4 N_NET12_20 0.00128722f
cc_56 N_C_4 N_NET12_3 0.00219243f
cc_57 N_MM2_g N_NET12_14 0.0353325f
cc_58 N_C_1 N_D_4 0.00108091f
cc_59 N_MM2_g N_MM3_g 0.00522093f
cc_60 N_C_4 N_D_4 0.00681636f
x_PM_OR4x2_ASAP7_75t_R%B VSS B N_MM6_g N_B_1 N_B_4 PM_OR4x2_ASAP7_75t_R%B
cc_61 N_MM6_g N_NET12_21 0.000210741f
cc_62 N_MM6_g N_NET12_4 0.00149219f
cc_63 N_MM6_g N_NET12_5 0.000344731f
cc_64 N_B_1 N_NET12_15 0.000711123f
cc_65 N_B_4 N_NET12_20 0.0011926f
cc_66 N_B_4 N_NET12_4 0.00232286f
cc_67 N_MM6_g N_NET12_15 0.0356501f
cc_68 N_B_1 N_C_1 0.00128681f
cc_69 N_MM6_g N_MM2_g 0.00542776f
cc_70 N_B_4 N_C_4 0.00761904f
x_PM_OR4x2_ASAP7_75t_R%NET12 VSS N_MM9_g N_MM9@2_g N_MM3_d N_MM2_d N_MM1_d
+ N_MM0_d N_MM7_d N_NET12_20 N_NET12_24 N_NET12_1 N_NET12_3 N_NET12_17
+ N_NET12_14 N_NET12_21 N_NET12_4 N_NET12_5 N_NET12_15 N_NET12_16 N_NET12_25
+ N_NET12_23 N_NET12_22 N_NET12_18 PM_OR4x2_ASAP7_75t_R%NET12
*END of OR4x2_ASAP7_75t_R.pxi
.ENDS
** Design:	OR5x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR5x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR5x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR5x1_ASAP7_75t_R%NET023 VSS 2 3 1
c1 1 VSS 0.000900038f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR5x1_ASAP7_75t_R%NET027 VSS 2 3 1
c1 1 VSS 0.000861049f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_OR5x1_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000867018f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_OR5x1_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000854785f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR5x1_ASAP7_75t_R%D VSS 10 3 1 4
c1 1 VSS 0.00392225f
c2 3 VSS 0.035438f
c3 4 VSS 0.00742644f
r1 10 9 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1360 $X2=0.2430 $Y2=0.1165
r2 4 9 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0935 $X2=0.2430 $Y2=0.1165
r3 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1355
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1360
+ $X2=0.2430 $Y2=0.1355
.ends

.subckt PM_OR5x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00441363f
.ends

.subckt PM_OR5x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00483246f
.ends

.subckt PM_OR5x1_ASAP7_75t_R%A VSS 11 3 1 4
c1 1 VSS 0.00510087f
c2 3 VSS 0.034839f
c3 4 VSS 0.00453338f
r1 11 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0810 $Y2=0.0985
r2 7 10 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1360 $X2=0.0915 $Y2=0.1360
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0905 $Y2=0.1360
r4 11 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1360
+ $X2=0.0810 $Y2=0.1360
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0810 $Y2=0.1360
r6 1 8 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0685 $Y2=0.1360
r7 3 6 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1360
r8 3 8 4.17867 $w=1.8386e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1360
r9 3 10 1.08747 $w=2.16729e-07 $l=1.05475e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1360
.ends

.subckt PM_OR5x1_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00428025f
c2 3 VSS 0.0352784f
c3 4 VSS 0.00725853f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1360 $X2=0.1890 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1360
+ $X2=0.1890 $Y2=0.1355
.ends

.subckt PM_OR5x1_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00346154f
c2 3 VSS 0.0348978f
c3 4 VSS 0.00685462f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1360
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_OR5x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00473964f
.ends

.subckt PM_OR5x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00458004f
.ends

.subckt PM_OR5x1_ASAP7_75t_R%E VSS 8 3 1 4
c1 1 VSS 0.00654559f
c2 3 VSS 0.0832594f
c3 4 VSS 0.00762114f
r1 8 4 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1360 $X2=0.2970 $Y2=0.1165
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1360
+ $X2=0.2970 $Y2=0.1355
.ends

.subckt PM_OR5x1_ASAP7_75t_R%NET024 VSS 15 54 55 58 59 63 68 16 26 4 3 21 19 20
+ 5 17 6 28 18 23 1 24 29
c1 1 VSS 0.00364552f
c2 3 VSS 0.00732642f
c3 4 VSS 0.00607878f
c4 5 VSS 0.00835585f
c5 6 VSS 0.00876097f
c6 15 VSS 0.0800026f
c7 16 VSS 0.00353752f
c8 17 VSS 0.00430243f
c9 18 VSS 0.0044151f
c10 19 VSS 0.00311281f
c11 20 VSS 0.00393805f
c12 21 VSS 0.0225616f
c13 22 VSS 0.00053728f
c14 23 VSS 0.00135467f
c15 24 VSS 0.00141329f
c16 25 VSS 0.00299406f
c17 26 VSS 0.00655307f
c18 27 VSS 0.00273291f
c19 28 VSS 0.000545266f
c20 29 VSS 0.00047742f
r1 68 67 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 19 67 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 4 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 64 65 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 26 61 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 26 64 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 63 62 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r8 16 62 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r9 60 61 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.2125
r10 20 25 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r11 20 60 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1350
r12 59 57 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r13 5 57 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r14 17 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r15 58 17 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r16 55 53 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2845 $Y2=0.0540
r17 6 53 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0540 $X2=0.2845 $Y2=0.0540
r18 18 6 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r19 54 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2555 $Y2=0.0540
r20 3 50 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r21 25 49 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r22 5 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r23 6 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r24 50 51 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0665 $Y2=0.0360
r25 49 50 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r26 48 51 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0710
+ $Y=0.0360 $X2=0.0665 $Y2=0.0360
r27 47 48 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0710 $Y2=0.0360
r28 46 47 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r29 45 46 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r30 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r31 42 43 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r32 42 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r33 41 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r34 40 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r35 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r36 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r37 21 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r38 21 39 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r39 27 38 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2835 $Y2=0.0360
r40 22 28 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0540 $X2=0.2970 $Y2=0.0665
r41 22 27 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0360
r42 23 29 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.0720 $X2=0.3510 $Y2=0.0720
r43 23 28 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.0720 $X2=0.2970 $Y2=0.0665
r44 29 35 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0935
r45 24 33 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1165 $X2=0.3510 $Y2=0.1360
r46 24 35 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1165 $X2=0.3510 $Y2=0.0935
r47 15 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1355
r48 1 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1355
+ $X2=0.3510 $Y2=0.1360
r49 4 19 1e-05
r50 3 16 1e-05
.ends

.subckt PM_OR5x1_ASAP7_75t_R%Y VSS 20 15 27 10 7 2 1 8 9 11
c1 1 VSS 0.00799623f
c2 2 VSS 0.00811983f
c3 7 VSS 0.00386434f
c4 8 VSS 0.00382569f
c5 9 VSS 0.00478609f
c6 10 VSS 0.00497016f
c7 11 VSS 0.00379667f
c8 12 VSS 0.0028682f
c9 13 VSS 0.00284658f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3760 $Y2=0.2025
r2 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r3 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r4 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r5 10 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r6 13 22 8.72783 $w=1.4982e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.4050 $Y2=0.1895
r7 13 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.2340 $X2=0.3915 $Y2=0.2340
r8 21 22 11.1348 $w=1.3e-08 $l=4.78e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1417 $X2=0.4050 $Y2=0.1895
r9 20 21 2.97317 $w=1.3e-08 $l=1.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1290 $X2=0.4050 $Y2=0.1417
r10 20 19 7.75356 $w=1.3e-08 $l=3.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1290 $X2=0.4050 $Y2=0.0957
r11 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0360
r12 11 19 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0540 $X2=0.4050 $Y2=0.0957
r13 12 17 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0360 $X2=0.3915 $Y2=0.0360
r14 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r15 9 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r16 1 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r17 7 1 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3760 $Y2=0.0675
r18 15 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
.ends


*
.SUBCKT OR5x1_ASAP7_75t_R VSS VDD A B C D E Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* E E
* Y Y
*
*

MM10 VSS N_MM10_g N_MM10_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 VSS N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 VSS N_MM8_g N_MM8_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 VSS N_MM6_g N_MM9_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 VSS N_MM11_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM10_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM2_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM7_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM8_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 VDD N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VDD N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR5x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR5x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR5x1_ASAP7_75t_R%NET023 VSS N_MM0_d N_MM4_s N_NET023_1
+ PM_OR5x1_ASAP7_75t_R%NET023
cc_1 N_NET023_1 N_MM10_g 0.0174959f
cc_2 N_NET023_1 N_MM2_g 0.0173895f
x_PM_OR5x1_ASAP7_75t_R%NET027 VSS N_MM6_s N_MM5_d N_NET027_1
+ PM_OR5x1_ASAP7_75t_R%NET027
cc_3 N_NET027_1 N_MM8_g 0.0175071f
cc_4 N_NET027_1 N_MM6_g 0.0173636f
x_PM_OR5x1_ASAP7_75t_R%NET29 VSS N_MM3_d N_MM5_s N_NET29_1
+ PM_OR5x1_ASAP7_75t_R%NET29
cc_5 N_NET29_1 N_MM7_g 0.0176318f
cc_6 N_NET29_1 N_MM8_g 0.0175084f
x_PM_OR5x1_ASAP7_75t_R%NET30 VSS N_MM4_d N_MM3_s N_NET30_1
+ PM_OR5x1_ASAP7_75t_R%NET30
cc_7 N_NET30_1 N_MM2_g 0.0176269f
cc_8 N_NET30_1 N_MM7_g 0.0175252f
x_PM_OR5x1_ASAP7_75t_R%D VSS D N_MM8_g N_D_1 N_D_4 PM_OR5x1_ASAP7_75t_R%D
cc_9 N_D_1 N_C_1 0.0017261f
cc_10 N_D_4 N_C_4 0.00677952f
cc_11 N_MM8_g N_MM7_g 0.00871804f
x_PM_OR5x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_OR5x1_ASAP7_75t_R%noxref_14
cc_12 N_noxref_14_1 N_MM10_g 0.00356505f
cc_13 N_noxref_14_1 N_NET024_3 0.00050372f
cc_14 N_noxref_14_1 N_NET024_16 0.0282766f
x_PM_OR5x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_OR5x1_ASAP7_75t_R%noxref_15
cc_15 N_noxref_15_1 N_MM10_g 0.00166313f
cc_16 N_noxref_15_1 N_NET024_4 0.00049938f
cc_17 N_noxref_15_1 N_NET024_19 0.0376257f
cc_18 N_noxref_15_1 N_noxref_14_1 0.0018934f
x_PM_OR5x1_ASAP7_75t_R%A VSS A N_MM10_g N_A_1 N_A_4 PM_OR5x1_ASAP7_75t_R%A
x_PM_OR5x1_ASAP7_75t_R%C VSS C N_MM7_g N_C_1 N_C_4 PM_OR5x1_ASAP7_75t_R%C
cc_19 N_C_1 N_B_1 0.00167659f
cc_20 N_C_4 N_B_4 0.00635516f
cc_21 N_MM7_g N_MM2_g 0.00876845f
x_PM_OR5x1_ASAP7_75t_R%B VSS B N_MM2_g N_B_1 N_B_4 PM_OR5x1_ASAP7_75t_R%B
cc_22 N_B_1 N_A_1 0.00146301f
cc_23 N_B_4 N_A_4 0.00558325f
cc_24 N_MM2_g N_MM10_g 0.00850017f
x_PM_OR5x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_OR5x1_ASAP7_75t_R%noxref_17
cc_25 N_noxref_17_1 N_MM11_g 0.00145317f
cc_26 N_noxref_17_1 N_Y_8 0.0384569f
cc_27 N_noxref_17_1 N_noxref_16_1 0.00177678f
x_PM_OR5x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_OR5x1_ASAP7_75t_R%noxref_16
cc_28 N_noxref_16_1 N_MM11_g 0.0014585f
cc_29 N_noxref_16_1 N_Y_7 0.0385868f
x_PM_OR5x1_ASAP7_75t_R%E VSS E N_MM6_g N_E_1 N_E_4 PM_OR5x1_ASAP7_75t_R%E
cc_30 N_E_1 N_D_1 0.00152928f
cc_31 N_E_4 N_D_4 0.00567693f
cc_32 N_MM6_g N_MM8_g 0.00849912f
x_PM_OR5x1_ASAP7_75t_R%NET024 VSS N_MM11_g N_MM8_s N_MM9_s N_MM2_s N_MM7_s
+ N_MM10_s N_MM0_s N_NET024_16 N_NET024_26 N_NET024_4 N_NET024_3 N_NET024_21
+ N_NET024_19 N_NET024_20 N_NET024_5 N_NET024_17 N_NET024_6 N_NET024_28
+ N_NET024_18 N_NET024_23 N_NET024_1 N_NET024_24 N_NET024_29
+ PM_OR5x1_ASAP7_75t_R%NET024
cc_33 N_NET024_16 N_MM10_g 0.011217f
cc_34 N_NET024_26 N_A_4 0.000571175f
cc_35 N_NET024_4 N_A_1 0.000698572f
cc_36 N_NET024_3 N_MM10_g 0.000749817f
cc_37 N_NET024_21 N_A_4 0.0012197f
cc_38 N_NET024_4 N_MM10_g 0.00194499f
cc_39 N_NET024_19 N_A_1 0.00198479f
cc_40 N_NET024_20 N_A_4 0.00853529f
cc_41 N_NET024_19 N_MM10_g 0.0497448f
cc_42 N_NET024_26 N_MM2_g 0.000202152f
cc_43 N_NET024_20 N_MM2_g 0.000216385f
cc_44 N_NET024_4 N_MM2_g 0.000350924f
cc_45 N_NET024_5 N_MM2_g 0.000709487f
cc_46 N_NET024_21 N_B_4 0.0012792f
cc_47 N_NET024_4 N_B_4 0.00214477f
cc_48 N_NET024_17 N_MM2_g 0.0262441f
cc_49 N_NET024_5 N_MM7_g 0.000710587f
cc_50 N_NET024_21 N_C_4 0.00128797f
cc_51 N_NET024_5 N_C_4 0.00179768f
cc_52 N_NET024_17 N_MM7_g 0.025883f
cc_53 N_NET024_6 N_MM8_g 0.000698158f
cc_54 N_NET024_21 N_D_4 0.00121109f
cc_55 N_NET024_28 N_D_4 0.0024982f
cc_56 N_NET024_18 N_MM8_g 0.0261183f
cc_57 N_NET024_23 N_MM6_g 0.000385406f
cc_58 N_NET024_6 N_MM6_g 0.000407112f
cc_59 N_NET024_28 N_MM6_g 0.000534994f
cc_60 N_NET024_1 N_E_1 0.00216731f
cc_61 N_NET024_24 N_E_4 0.00363987f
cc_62 N_NET024_18 N_MM6_g 0.0109287f
cc_63 N_MM11_g N_MM6_g 0.017498f
x_PM_OR5x1_ASAP7_75t_R%Y VSS Y N_MM1_s N_MM11_s N_Y_10 N_Y_7 N_Y_2 N_Y_1 N_Y_8
+ N_Y_9 N_Y_11 PM_OR5x1_ASAP7_75t_R%Y
cc_64 N_Y_10 N_E_4 0.00196772f
cc_65 N_Y_7 N_NET024_29 0.000180589f
cc_66 N_Y_7 N_NET024_23 0.000456262f
cc_67 N_Y_2 N_NET024_1 0.000850689f
cc_68 N_Y_2 N_MM11_g 0.00105953f
cc_69 N_Y_1 N_MM11_g 0.00139203f
cc_70 N_Y_8 N_NET024_1 0.0015691f
cc_71 N_Y_9 N_NET024_29 0.00241713f
cc_72 N_Y_11 N_NET024_24 0.00468232f
cc_73 N_Y_8 N_MM11_g 0.0152198f
cc_74 N_Y_7 N_MM11_g 0.0551357f
*END of OR5x1_ASAP7_75t_R.pxi
.ENDS
** Design:	OR5x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "OR5x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "OR5x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_OR5x2_ASAP7_75t_R%NET027 VSS 2 3 1
c1 1 VSS 0.000890568f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2700 $Y2=0.2025
.ends

.subckt PM_OR5x2_ASAP7_75t_R%NET29 VSS 2 3 1
c1 1 VSS 0.000869499f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_OR5x2_ASAP7_75t_R%NET30 VSS 2 3 1
c1 1 VSS 0.000842815f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_OR5x2_ASAP7_75t_R%NET023 VSS 2 3 1
c1 1 VSS 0.000902512f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_OR5x2_ASAP7_75t_R%A VSS 11 3 1 4
c1 1 VSS 0.00524617f
c2 3 VSS 0.034912f
c3 4 VSS 0.00457955f
r1 11 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0810 $Y2=0.0985
r2 7 10 0.966062 $w=1.465e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0905
+ $Y=0.1360 $X2=0.0915 $Y2=0.1360
r3 6 7 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1360 $X2=0.0905 $Y2=0.1360
r4 11 6 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1360
+ $X2=0.0810 $Y2=0.1360
r5 1 6 3.67195 $w=1.8e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0810 $Y2=0.1360
r6 1 8 4.05727 $w=1.24167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1360 $X2=0.0685 $Y2=0.1360
r7 3 6 3.79335 $w=1.28e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1360
r8 3 8 4.17867 $w=1.8386e-07 $l=1.25399e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1360
r9 3 10 1.08747 $w=2.16729e-07 $l=1.05475e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0915 $Y2=0.1360
.ends

.subckt PM_OR5x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0423818f
.ends

.subckt PM_OR5x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0423821f
.ends

.subckt PM_OR5x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00442797f
.ends

.subckt PM_OR5x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00483593f
.ends

.subckt PM_OR5x2_ASAP7_75t_R%E VSS 8 3 4 1
c1 1 VSS 0.00669667f
c2 3 VSS 0.0834378f
c3 4 VSS 0.00890837f
r1 8 4 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1360 $X2=0.2970 $Y2=0.1165
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1360
+ $X2=0.2970 $Y2=0.1355
.ends

.subckt PM_OR5x2_ASAP7_75t_R%B VSS 8 3 1 4
c1 1 VSS 0.00367676f
c2 3 VSS 0.0350081f
c3 4 VSS 0.00692817f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1360 $X2=0.1350 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1360
+ $X2=0.1350 $Y2=0.1355
.ends

.subckt PM_OR5x2_ASAP7_75t_R%C VSS 8 3 1 4
c1 1 VSS 0.00406711f
c2 3 VSS 0.0352217f
c3 4 VSS 0.00733586f
r1 8 4 8.74462 $w=1.3e-08 $l=3.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1360 $X2=0.1890 $Y2=0.0985
r2 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1355
r3 8 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1360
+ $X2=0.1890 $Y2=0.1355
.ends

.subckt PM_OR5x2_ASAP7_75t_R%D VSS 10 3 1 4
c1 1 VSS 0.00411577f
c2 3 VSS 0.0355142f
c3 4 VSS 0.00736146f
r1 10 9 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1360 $X2=0.2430 $Y2=0.1165
r2 4 9 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0935 $X2=0.2430 $Y2=0.1165
r3 3 1 3.81699 $w=1.23e-07 $l=5e-10 $layer=LIG $thickness=5.2e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1355
r4 10 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1360
+ $X2=0.2430 $Y2=0.1355
.ends

.subckt PM_OR5x2_ASAP7_75t_R%Y VSS 23 16 17 30 31 7 11 1 2 9 8
c1 1 VSS 0.0102042f
c2 2 VSS 0.0116214f
c3 7 VSS 0.00463308f
c4 8 VSS 0.00454934f
c5 9 VSS 0.011f
c6 10 VSS 0.00972395f
c7 11 VSS 0.00766542f
c8 12 VSS 0.00336496f
c9 13 VSS 0.0034551f
r1 31 29 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 2 29 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 30 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r6 26 27 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r7 10 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r8 13 25 8.72783 $w=1.4982e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4590 $Y2=0.1895
r9 13 27 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4185 $Y2=0.2340
r10 24 25 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1510 $X2=0.4590 $Y2=0.1895
r11 23 24 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1510
r12 23 22 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1050
r13 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r14 11 22 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.1050
r15 12 21 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4185 $Y2=0.0360
r16 20 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r17 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r18 9 19 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3620
+ $Y=0.0360 $X2=0.3665 $Y2=0.0360
r19 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r20 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r21 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r22 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r23 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
.ends

.subckt PM_OR5x2_ASAP7_75t_R%NET024 VSS 15 16 63 64 67 68 72 77 17 27 4 3 22 20
+ 21 5 18 6 29 19 24 1 25 30
c1 1 VSS 0.00752739f
c2 3 VSS 0.00750828f
c3 4 VSS 0.00626572f
c4 5 VSS 0.00836538f
c5 6 VSS 0.0087727f
c6 15 VSS 0.0804021f
c7 16 VSS 0.0808426f
c8 17 VSS 0.00440554f
c9 18 VSS 0.00514715f
c10 19 VSS 0.00526709f
c11 20 VSS 0.00427123f
c12 21 VSS 0.00615767f
c13 22 VSS 0.0230614f
c14 23 VSS 0.000525413f
c15 24 VSS 0.00139708f
c16 25 VSS 0.00221435f
c17 26 VSS 0.00329981f
c18 27 VSS 0.00713749f
c19 28 VSS 0.00270352f
c20 29 VSS 0.000543233f
c21 30 VSS 0.000506555f
r1 77 76 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 20 76 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 4 74 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 73 74 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 27 70 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 27 73 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 72 71 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r8 17 71 0.231482 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0540 $X2=0.0685 $Y2=0.0540
r9 69 70 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.2125
r10 21 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0575 $X2=0.0270 $Y2=0.0360
r11 21 69 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0575 $X2=0.0270 $Y2=0.1350
r12 68 66 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r13 5 66 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1620 $Y=0.0540 $X2=0.1765 $Y2=0.0540
r14 18 5 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0540 $X2=0.1620 $Y2=0.0540
r15 67 18 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0540 $X2=0.1475 $Y2=0.0540
r16 64 62 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0540 $X2=0.2845 $Y2=0.0540
r17 6 62 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0540 $X2=0.2845 $Y2=0.0540
r18 19 6 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0540 $X2=0.2700 $Y2=0.0540
r19 63 19 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0540 $X2=0.2555 $Y2=0.0540
r20 3 59 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0540
+ $X2=0.0540 $Y2=0.0360
r21 26 58 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r22 5 52 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1620 $Y=0.0540
+ $X2=0.1620 $Y2=0.0360
r23 6 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r24 59 60 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.0665 $Y2=0.0360
r25 58 59 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r26 57 60 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0710
+ $Y=0.0360 $X2=0.0665 $Y2=0.0360
r27 56 57 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.0710 $Y2=0.0360
r28 55 56 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r29 54 55 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r30 52 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r31 51 52 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r32 51 54 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1485
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r33 50 53 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0360 $X2=0.1755 $Y2=0.0360
r34 49 50 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1890 $Y2=0.0360
r35 48 49 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r36 46 47 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.2835 $Y2=0.0360
r37 22 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r38 22 48 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.0360 $X2=0.2430 $Y2=0.0360
r39 28 47 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0360 $X2=0.2835 $Y2=0.0360
r40 23 29 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2970 $Y=0.0540 $X2=0.2970 $Y2=0.0665
r41 23 28 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0540 $X2=0.2970 $Y2=0.0360
r42 24 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.0720 $X2=0.3510 $Y2=0.0720
r43 24 29 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.0720 $X2=0.2970 $Y2=0.0665
r44 30 43 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0935
r45 16 39 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r46 25 41 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1165 $X2=0.3510 $Y2=0.1360
r47 25 43 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1165 $X2=0.3510 $Y2=0.0935
r48 37 39 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r49 36 37 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3780 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r50 35 36 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3780 $Y2=0.1350
r51 33 35 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3605 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r52 32 33 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3605 $Y2=0.1350
r53 32 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1360
r54 1 32 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r55 1 34 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3405 $Y2=0.1350
r56 15 32 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r57 15 34 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r58 15 35 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r59 4 20 1e-05
r60 3 17 1e-05
.ends


*
.SUBCKT OR5x2_ASAP7_75t_R VSS VDD A B C D E Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* D D
* E E
* Y Y
*
*

MM10 VSS N_MM10_g N_MM10_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM2 VSS N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM7 VSS N_MM7_g N_MM7_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM8 VSS N_MM5_g N_MM8_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM9 VSS N_MM6_g N_MM9_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 VSS N_MM11_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1@2 VSS N_MM11@2_g N_MM1@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM10_g N_MM0_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM2_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM7_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 VDD N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VDD N_MM11_g N_MM11_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 VDD N_MM11@2_g N_MM11@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "OR5x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "OR5x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_OR5x2_ASAP7_75t_R%NET027 VSS N_MM5_d N_MM6_s N_NET027_1
+ PM_OR5x2_ASAP7_75t_R%NET027
cc_1 N_NET027_1 N_MM5_g 0.0174919f
cc_2 N_NET027_1 N_MM6_g 0.0173493f
x_PM_OR5x2_ASAP7_75t_R%NET29 VSS N_MM5_s N_MM3_d N_NET29_1
+ PM_OR5x2_ASAP7_75t_R%NET29
cc_3 N_NET29_1 N_MM7_g 0.0176348f
cc_4 N_NET29_1 N_MM5_g 0.0175028f
x_PM_OR5x2_ASAP7_75t_R%NET30 VSS N_MM4_d N_MM3_s N_NET30_1
+ PM_OR5x2_ASAP7_75t_R%NET30
cc_5 N_NET30_1 N_MM2_g 0.0176305f
cc_6 N_NET30_1 N_MM7_g 0.0175335f
x_PM_OR5x2_ASAP7_75t_R%NET023 VSS N_MM0_d N_MM4_s N_NET023_1
+ PM_OR5x2_ASAP7_75t_R%NET023
cc_7 N_NET023_1 N_MM10_g 0.0174942f
cc_8 N_NET023_1 N_MM2_g 0.0173888f
x_PM_OR5x2_ASAP7_75t_R%A VSS A N_MM10_g N_A_1 N_A_4 PM_OR5x2_ASAP7_75t_R%A
x_PM_OR5x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_OR5x2_ASAP7_75t_R%noxref_16
cc_9 N_noxref_16_1 N_MM11@2_g 0.00146947f
cc_10 N_noxref_16_1 N_Y_7 0.000853276f
x_PM_OR5x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_OR5x2_ASAP7_75t_R%noxref_17
cc_11 N_noxref_17_1 N_MM11@2_g 0.00147484f
cc_12 N_noxref_17_1 N_Y_8 0.000855051f
cc_13 N_noxref_17_1 N_noxref_16_1 0.00177287f
x_PM_OR5x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_OR5x2_ASAP7_75t_R%noxref_14
cc_14 N_noxref_14_1 N_MM10_g 0.00357957f
cc_15 N_noxref_14_1 N_NET024_21 0.000362142f
cc_16 N_noxref_14_1 N_NET024_3 0.00050372f
cc_17 N_noxref_14_1 N_NET024_17 0.0279142f
x_PM_OR5x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_OR5x2_ASAP7_75t_R%noxref_15
cc_18 N_noxref_15_1 N_MM10_g 0.00166311f
cc_19 N_noxref_15_1 N_NET024_4 0.00049645f
cc_20 N_noxref_15_1 N_NET024_20 0.0376101f
cc_21 N_noxref_15_1 N_noxref_14_1 0.00189248f
x_PM_OR5x2_ASAP7_75t_R%E VSS E N_MM6_g N_E_4 N_E_1 PM_OR5x2_ASAP7_75t_R%E
cc_22 N_MM6_g N_D_1 0.00156233f
cc_23 N_E_4 N_D_4 0.00561556f
cc_24 N_MM6_g N_MM5_g 0.00831754f
x_PM_OR5x2_ASAP7_75t_R%B VSS B N_MM2_g N_B_1 N_B_4 PM_OR5x2_ASAP7_75t_R%B
cc_25 N_B_1 N_A_1 0.00146301f
cc_26 N_B_4 N_A_4 0.00557948f
cc_27 N_MM2_g N_MM10_g 0.00850017f
x_PM_OR5x2_ASAP7_75t_R%C VSS C N_MM7_g N_C_1 N_C_4 PM_OR5x2_ASAP7_75t_R%C
cc_28 N_C_1 N_B_1 0.00156042f
cc_29 N_C_4 N_B_4 0.0066212f
cc_30 N_MM7_g N_MM2_g 0.00876845f
x_PM_OR5x2_ASAP7_75t_R%D VSS D N_MM5_g N_D_1 N_D_4 PM_OR5x2_ASAP7_75t_R%D
cc_31 N_D_1 N_C_1 0.00160977f
cc_32 N_D_4 N_C_4 0.00672511f
cc_33 N_MM5_g N_MM7_g 0.00872153f
x_PM_OR5x2_ASAP7_75t_R%Y VSS Y N_MM1_s N_MM1@2_s N_MM11_s N_MM11@2_s N_Y_7
+ N_Y_11 N_Y_1 N_Y_2 N_Y_9 N_Y_8 PM_OR5x2_ASAP7_75t_R%Y
cc_34 N_Y_7 N_NET024_30 0.000232877f
cc_35 N_Y_7 N_NET024_25 0.000307148f
cc_36 N_Y_7 N_NET024_24 0.000531549f
cc_37 N_Y_7 N_NET024_1 0.000532107f
cc_38 N_Y_11 N_NET024_1 0.000936227f
cc_39 N_Y_1 N_NET024_25 0.00148262f
cc_40 N_Y_2 N_MM11_g 0.00203422f
cc_41 N_Y_1 N_MM11_g 0.00234603f
cc_42 N_Y_9 N_NET024_30 0.00299448f
cc_43 N_Y_8 N_NET024_1 0.00455275f
cc_44 N_Y_8 N_MM11_g 0.0300419f
cc_45 N_Y_7 N_MM11@2_g 0.0373051f
cc_46 N_Y_7 N_MM11_g 0.0697629f
x_PM_OR5x2_ASAP7_75t_R%NET024 VSS N_MM11_g N_MM11@2_g N_MM8_s N_MM9_s N_MM2_s
+ N_MM7_s N_MM10_s N_MM0_s N_NET024_17 N_NET024_27 N_NET024_4 N_NET024_3
+ N_NET024_22 N_NET024_20 N_NET024_21 N_NET024_5 N_NET024_18 N_NET024_6
+ N_NET024_29 N_NET024_19 N_NET024_24 N_NET024_1 N_NET024_25 N_NET024_30
+ PM_OR5x2_ASAP7_75t_R%NET024
cc_47 N_NET024_17 N_MM10_g 0.011217f
cc_48 N_NET024_27 N_A_4 0.000540932f
cc_49 N_NET024_4 N_A_1 0.000698572f
cc_50 N_NET024_3 N_MM10_g 0.000749817f
cc_51 N_NET024_22 N_A_4 0.00105001f
cc_52 N_NET024_4 N_MM10_g 0.00194546f
cc_53 N_NET024_20 N_A_1 0.00198479f
cc_54 N_NET024_21 N_A_4 0.00859496f
cc_55 N_NET024_20 N_MM10_g 0.0497322f
cc_56 N_NET024_21 N_MM2_g 0.000193133f
cc_57 N_NET024_27 N_MM2_g 0.00020436f
cc_58 N_NET024_4 N_MM2_g 0.000348453f
cc_59 N_NET024_5 N_MM2_g 0.000709487f
cc_60 N_NET024_22 N_B_4 0.00112928f
cc_61 N_NET024_4 N_B_4 0.00218499f
cc_62 N_NET024_18 N_MM2_g 0.0262819f
cc_63 N_NET024_5 N_MM7_g 0.000710587f
cc_64 N_NET024_22 N_C_4 0.00110325f
cc_65 N_NET024_5 N_C_4 0.00177259f
cc_66 N_NET024_18 N_MM7_g 0.0258003f
cc_67 N_NET024_6 N_MM5_g 0.00084037f
cc_68 N_NET024_22 N_D_4 0.00106042f
cc_69 N_NET024_29 N_D_4 0.0026937f
cc_70 N_NET024_19 N_MM5_g 0.0259918f
cc_71 N_NET024_24 N_MM6_g 0.000379516f
cc_72 N_NET024_6 N_MM6_g 0.000420168f
cc_73 N_NET024_29 N_MM6_g 0.00056909f
cc_74 N_NET024_1 N_E_1 0.00200808f
cc_75 N_NET024_25 N_E_4 0.00364083f
cc_76 N_NET024_19 N_MM6_g 0.0109297f
cc_77 N_MM11_g N_MM6_g 0.0174986f
*END of OR5x2_ASAP7_75t_R.pxi
.ENDS
** Design:	XOR2x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XOR2x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XOR2x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XOR2x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.042214f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0422992f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%NET047 VSS 2 3 1
c1 1 VSS 0.00103441f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5400 $Y2=0.0675
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%NET048 VSS 2 3 1
c1 1 VSS 0.000993129f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00654585f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%NET047__2 VSS 2 3 1
c1 1 VSS 0.00102628f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0420734f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00631483f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00617239f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0048035f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00603065f
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%NET019 VSS 19 41 42 45 46 48 14 2 17 15 1 3 13 16
+ 4
c1 1 VSS 0.00699321f
c2 2 VSS 0.00702988f
c3 3 VSS 0.00711838f
c4 4 VSS 0.00804985f
c5 13 VSS 0.00371783f
c6 14 VSS 0.00333708f
c7 15 VSS 0.00332985f
c8 16 VSS 0.00343391f
c9 17 VSS 0.033465f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r2 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r3 46 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r4 3 44 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r5 15 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r6 45 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r7 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r8 2 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r9 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r10 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r11 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r12 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r13 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r14 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r15 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.2340 $X2=0.5805 $Y2=0.2340
r16 34 35 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5420
+ $Y=0.2340 $X2=0.5670 $Y2=0.2340
r17 33 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5240
+ $Y=0.2340 $X2=0.5420 $Y2=0.2340
r18 32 33 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5240 $Y2=0.2340
r19 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.2340 $X2=0.5130 $Y2=0.2340
r20 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4995 $Y2=0.2340
r21 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r22 28 29 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4430
+ $Y=0.2340 $X2=0.4725 $Y2=0.2340
r23 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.4430 $Y2=0.2340
r24 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r25 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.2340 $X2=0.4050 $Y2=0.2340
r26 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.2340 $X2=0.3915 $Y2=0.2340
r27 23 24 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r28 22 23 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3440
+ $Y=0.2340 $X2=0.3670 $Y2=0.2340
r29 21 22 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3010
+ $Y=0.2340 $X2=0.3440 $Y2=0.2340
r30 20 21 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3010 $Y2=0.2340
r31 17 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r32 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r33 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r34 13 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r35 1 13 1e-05
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%Y VSS 32 23 45 46 51 54 55 18 19 4 16 14 13 1 20
+ 15 17 2 3
c1 1 VSS 0.00592524f
c2 2 VSS 0.00954605f
c3 3 VSS 0.00286554f
c4 4 VSS 0.00620528f
c5 13 VSS 0.00308504f
c6 14 VSS 0.00441854f
c7 15 VSS 0.00261048f
c8 16 VSS 0.00203108f
c9 17 VSS 0.0172999f
c10 18 VSS 0.00168838f
c11 19 VSS 0.0137298f
c12 20 VSS 0.000268981f
c13 21 VSS 0.00206796f
r1 55 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r2 3 53 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r3 16 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r4 54 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 15 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r6 51 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r7 3 48 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.1840
r8 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0360
r9 48 49 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.1840 $X2=0.4455 $Y2=0.1840
r10 20 35 3.94987 $w=1.50455e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1840 $X2=0.4590 $Y2=0.1620
r11 20 49 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1840 $X2=0.4455 $Y2=0.1840
r12 46 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r13 2 44 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r14 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r15 45 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r16 39 40 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r17 38 39 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5510
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r18 37 38 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5240
+ $Y=0.0360 $X2=0.5510 $Y2=0.0360
r19 36 37 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5240 $Y2=0.0360
r20 19 21 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r21 19 36 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r22 34 35 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1335 $X2=0.4590 $Y2=0.1620
r23 33 34 6.58761 $w=1.3e-08 $l=2.83e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1052 $X2=0.4590 $Y2=0.1335
r24 32 33 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0920 $X2=0.4590 $Y2=0.1052
r25 32 31 1.34084 $w=1.3e-08 $l=5.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0920 $X2=0.4590 $Y2=0.0862
r26 30 31 3.32295 $w=1.3e-08 $l=1.42e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0720 $X2=0.4590 $Y2=0.0862
r27 18 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r28 18 30 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0720
r29 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r30 21 29 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r31 28 29 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r32 27 28 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r33 26 27 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.0360 $X2=0.4205 $Y2=0.0360
r34 25 26 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3465
+ $Y=0.0360 $X2=0.4160 $Y2=0.0360
r35 24 25 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3465 $Y2=0.0360
r36 17 24 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r37 1 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r38 23 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r39 13 22 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r40 1 13 1e-05
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%NET036 VSS 9 10 48 51 52 11 15 1 4 17 13 3 16 12
+ 19 20
c1 1 VSS 0.00581291f
c2 3 VSS 0.0123178f
c3 4 VSS 0.00793939f
c4 9 VSS 0.0434559f
c5 10 VSS 0.0435338f
c6 11 VSS 0.00779618f
c7 12 VSS 0.00540202f
c8 13 VSS 0.00960716f
c9 14 VSS 0.00167946f
c10 15 VSS 0.00236814f
c11 16 VSS 0.00480741f
c12 17 VSS 0.00163302f
c13 18 VSS 0.00359067f
c14 19 VSS 0.00145703f
c15 20 VSS 0.00130759f
r1 52 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r2 3 50 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r3 11 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r4 51 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r5 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1120 $Y2=0.0360
r6 12 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r7 48 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r8 43 44 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r9 13 18 3.94193 $w=1.70327e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1590 $Y=0.0360 $X2=0.1835 $Y2=0.0360
r10 13 44 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r11 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1750 $Y=0.2025
+ $X2=0.1830 $Y2=0.1740
r12 39 40 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1570 $X2=0.1830 $Y2=0.1740
r13 38 39 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1375 $X2=0.1830 $Y2=0.1570
r14 15 19 6.19173 $w=1.44844e-08 $l=3.1504e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1830 $Y=0.1035 $X2=0.1835 $Y2=0.0720
r15 15 38 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1035 $X2=0.1830 $Y2=0.1375
r16 14 19 2.64331 $w=1.65e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.0540 $X2=0.1835 $Y2=0.0720
r17 14 18 2.23928 $w=1.65e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.0540 $X2=0.1835 $Y2=0.0360
r18 19 37 3.27685 $w=1.54359e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1835 $Y=0.0720 $X2=0.2030 $Y2=0.0720
r19 36 37 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2345
+ $Y=0.0720 $X2=0.2030 $Y2=0.0720
r20 35 36 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2805
+ $Y=0.0720 $X2=0.2345 $Y2=0.0720
r21 34 35 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3350
+ $Y=0.0720 $X2=0.2805 $Y2=0.0720
r22 16 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3805 $Y=0.0720 $X2=0.4050 $Y2=0.0720
r23 16 34 10.6101 $w=1.3e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3805
+ $Y=0.0720 $X2=0.3350 $Y2=0.0720
r24 20 31 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0720 $X2=0.4050 $Y2=0.1035
r25 10 29 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r26 17 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r27 17 31 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1035
r28 27 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r29 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r30 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r31 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r32 22 23 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4145 $Y2=0.1350
r33 1 22 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r34 1 24 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.3945 $Y2=0.1350
r35 9 22 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r36 9 24 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r37 9 25 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%B VSS 37 5 6 7 9 1 8 10 11 2 12
c1 1 VSS 0.00705329f
c2 2 VSS 0.0026197f
c3 5 VSS 0.0436342f
c4 6 VSS 0.0435062f
c5 7 VSS 0.0431214f
c6 8 VSS 0.00291279f
c7 9 VSS 0.00477527f
c8 10 VSS 0.00101425f
c9 11 VSS 0.00130417f
c10 12 VSS 0.0388181f
r1 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r2 7 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 11 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0720 $X2=0.5670
+ $Y2=0.0810
r4 44 45 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1220 $X2=0.5670 $Y2=0.1350
r5 43 44 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1040 $X2=0.5670 $Y2=0.1220
r6 9 43 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0855 $X2=0.5670 $Y2=0.1040
r7 9 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.0855 $X2=0.5670
+ $Y2=0.0810
r8 9 11 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0855 $X2=0.5670 $Y2=0.0720
r9 40 41 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.5425
+ $Y=0.0810 $X2=0.5670 $Y2=0.0810
r10 39 40 30.3147 $w=1.3e-08 $l=1.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.4125
+ $Y=0.0810 $X2=0.5425 $Y2=0.0810
r11 38 39 36.3193 $w=1.3e-08 $l=1.558e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2567 $Y=0.0810 $X2=0.4125 $Y2=0.0810
r12 37 38 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M2 $thickness=3.6e-08 $X=0.2150
+ $Y=0.0810 $X2=0.2567 $Y2=0.0810
r13 37 36 8.33653 $w=1.3e-08 $l=3.58e-08 $layer=M2 $thickness=3.6e-08 $X=0.2150
+ $Y=0.0810 $X2=0.1792 $Y2=0.0810
r14 35 36 10.3186 $w=1.3e-08 $l=4.42e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0810 $X2=0.1792 $Y2=0.0810
r15 12 35 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1235
+ $Y=0.0810 $X2=0.1350 $Y2=0.0810
r16 10 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.0855
r17 10 35 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.0720 $X2=0.1350
+ $Y2=0.0810
r18 31 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0855 $X2=0.1350 $Y2=0.1080
r19 31 35 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.0855 $X2=0.1350
+ $Y2=0.0810
r20 8 29 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1350
r21 8 32 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1080
r22 5 24 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r23 24 25 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r24 24 29 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r25 21 25 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1445 $Y2=0.1350
r26 20 21 38.4626 $w=9.3e-09 $l=1.65e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1640 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r27 19 20 58.2767 $w=9.3e-09 $l=2.5e-08 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r28 18 19 93.2428 $w=9.3e-09 $l=4e-08 $layer=LIG $thickness=4.8e-08 $X=0.2290
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r29 17 18 95.5738 $w=9.3e-09 $l=4.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2290 $Y2=0.1350
r30 16 17 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r31 6 1 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r32 1 27 7.05813 $w=1.53909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3080 $Y2=0.1350
r33 6 16 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r34 6 27 2.64573 $w=2.07209e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3080 $Y2=0.1350
.ends

.subckt PM_XOR2x1_ASAP7_75t_R%A VSS 34 7 8 9 18 2 11 1 16 12 17 23 10 15 13 3
+ 25 21 14 22 24
c1 1 VSS 0.00882232f
c2 2 VSS 0.0039195f
c3 3 VSS 0.0042635f
c4 7 VSS 0.0818714f
c5 8 VSS 0.0815403f
c6 9 VSS 0.0814524f
c7 10 VSS 0.0120573f
c8 11 VSS 0.00854454f
c9 12 VSS 0.0021412f
c10 13 VSS 0.0205157f
c11 14 VSS 0.000361735f
c12 15 VSS 0.000904674f
c13 16 VSS 0.00105767f
c14 17 VSS 0.000401638f
c15 18 VSS 0.00234151f
c16 19 VSS 0.00200924f
c17 20 VSS 0.00488933f
c18 21 VSS 0.000252867f
c19 22 VSS 0.00285162f
c20 23 VSS 0.000234423f
c21 24 VSS 0.000639902f
c22 25 VSS 0.0140191f
r1 2 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r2 8 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 3 63 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r4 9 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 17 67 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3325
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 17 23 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3325 $Y=0.1350 $X2=0.3140 $Y2=0.1350
r7 63 64 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1465
r8 61 64 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1620 $X2=0.5130 $Y2=0.1465
r9 18 60 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1775 $X2=0.5130 $Y2=0.1865
r10 18 61 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1775 $X2=0.5130 $Y2=0.1620
r11 23 55 1.03257 $w=2.06696e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3140 $Y=0.1350 $X2=0.3140 $Y2=0.1465
r12 58 60 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.1890
+ $X2=0.5130 $Y2=0.1865
r13 57 58 23.2024 $w=1.3e-08 $l=9.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.4135
+ $Y=0.1890 $X2=0.5130 $Y2=0.1890
r14 56 57 23.2024 $w=1.3e-08 $l=9.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1890 $X2=0.4135 $Y2=0.1890
r15 25 56 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.3015
+ $Y=0.1890 $X2=0.3140 $Y2=0.1890
r16 54 55 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1620 $X2=0.3140 $Y2=0.1465
r17 53 56 70.3248 $w=5e-09 $l=1.8e-08 $layer=V1 $X=0.3140 $Y=0.1825 $X2=0.3140
+ $Y2=0.1890
r18 16 53 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1775 $X2=0.3140 $Y2=0.1825
r19 16 54 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1775 $X2=0.3140 $Y2=0.1620
r20 51 52 0.255111 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1990 $X2=0.3140 $Y2=0.2015
r21 50 51 0.357156 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1955 $X2=0.3140 $Y2=0.1990
r22 24 49 6.12133 $w=1.37018e-08 $l=3.38711e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3140 $Y=0.1890 $X2=0.2805 $Y2=0.1940
r23 24 50 0.663289 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1890 $X2=0.3140 $Y2=0.1955
r24 24 53 0.991152 $w=1.60769e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3140 $Y=0.1890 $X2=0.3140 $Y2=0.1825
r25 24 56 27.048 $w=1.3e-08 $l=1.8e-08 $layer=V1 $X=0.3140 $Y=0.1890 $X2=0.3140
+ $Y2=0.1890
r26 49 50 5.96826 $w=1.3463e-08 $l=3.35336e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2805 $Y=0.1940 $X2=0.3140 $Y2=0.1955
r27 49 52 5.86622 $w=1.32885e-08 $l=3.43293e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2805 $Y=0.1940 $X2=0.3140 $Y2=0.2015
r28 15 21 3.68021 $w=1.4875e-08 $l=2.15523e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2435 $Y=0.1940 $X2=0.2220 $Y2=0.1955
r29 15 49 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2435
+ $Y=0.1940 $X2=0.2805 $Y2=0.1940
r30 14 22 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2220
+ $Y=0.2140 $X2=0.2220 $Y2=0.2340
r31 14 21 3.33042 $w=1.5027e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2220 $Y=0.2140 $X2=0.2220 $Y2=0.1955
r32 22 47 2.89809 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2220 $Y=0.2340 $X2=0.2025 $Y2=0.2340
r33 46 47 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.2340 $X2=0.2025 $Y2=0.2340
r34 45 46 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.2340 $X2=0.1830 $Y2=0.2340
r35 44 45 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1590 $Y2=0.2340
r36 43 44 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1165
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r37 42 43 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0995
+ $Y=0.2340 $X2=0.1165 $Y2=0.2340
r38 41 42 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0850
+ $Y=0.2340 $X2=0.0995 $Y2=0.2340
r39 13 20 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.2340 $X2=0.0270 $Y2=0.2340
r40 13 41 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.2340 $X2=0.0850 $Y2=0.2340
r41 20 40 4.76361 $w=1.62073e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2065
r42 39 40 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1685 $X2=0.0270 $Y2=0.2065
r43 11 19 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1465 $X2=0.0270 $Y2=0.1350
r44 11 39 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1465 $X2=0.0270 $Y2=0.1685
r45 10 19 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r46 34 12 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r47 12 19 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r48 34 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r49 30 32 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r50 1 29 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r51 1 30 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r52 7 29 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r53 7 30 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends


*
.SUBCKT XOR2x1_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM0 VSS N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM5_g N_MM10@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 VSS N_MM4_g N_MM11@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 VSS N_MM6_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 VSS N_MM6@2_g N_MM9@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VSS N_MM4@2_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM5@2_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM0_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM1_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 VDD N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 VDD N_MM4_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM6@2_g N_MM6@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 VDD N_MM4@2_g N_MM4@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 VDD N_MM5@2_g N_MM5@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XOR2x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XOR2x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XOR2x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_A_1 0.000239215f
cc_2 N_noxref_12_1 N_MM0_g 0.00229937f
cc_3 N_noxref_12_1 N_noxref_11_1 0.00174589f
x_PM_XOR2x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_11
cc_4 N_noxref_11_1 N_A_1 0.000238356f
cc_5 N_noxref_11_1 N_MM0_g 0.00222976f
x_PM_XOR2x1_ASAP7_75t_R%NET047 VSS N_MM11_s N_MM10_d N_NET047_1
+ PM_XOR2x1_ASAP7_75t_R%NET047
cc_6 N_NET047_1 N_MM4@2_g 0.0174109f
cc_7 N_NET047_1 N_MM5@2_g 0.0173553f
x_PM_XOR2x1_ASAP7_75t_R%NET048 VSS N_MM3_s N_MM2_d N_NET048_1
+ PM_XOR2x1_ASAP7_75t_R%NET048
cc_8 N_NET048_1 N_MM0_g 0.0173137f
cc_9 N_NET048_1 N_MM1_g 0.0172255f
x_PM_XOR2x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_15
cc_10 N_noxref_15_1 N_B_1 0.00112832f
cc_11 N_noxref_15_1 N_MM5_g 0.00234367f
cc_12 N_noxref_15_1 N_Y_13 0.0355f
cc_13 N_noxref_15_1 N_noxref_13_1 0.00745617f
x_PM_XOR2x1_ASAP7_75t_R%NET047__2 VSS N_MM10@2_d N_MM11@2_s N_NET047__2_1
+ PM_XOR2x1_ASAP7_75t_R%NET047__2
cc_14 N_NET047__2_1 N_MM4_g 0.0172275f
cc_15 N_NET047__2_1 N_MM5_g 0.0173927f
x_PM_XOR2x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_13
cc_16 N_noxref_13_1 N_B_1 0.00111923f
cc_17 N_noxref_13_1 N_MM1_g 0.00232431f
x_PM_XOR2x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_18
cc_18 N_noxref_18_1 N_MM5@2_g 0.00163765f
cc_19 N_noxref_18_1 N_NET019_16 0.0360971f
cc_20 N_noxref_18_1 N_Y_15 0.000551921f
cc_21 N_noxref_18_1 N_noxref_17_1 0.00179021f
x_PM_XOR2x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_17
cc_22 N_noxref_17_1 N_MM5@2_g 0.00170615f
cc_23 N_noxref_17_1 N_NET019_16 0.000561219f
cc_24 N_noxref_17_1 N_Y_15 0.0362398f
x_PM_XOR2x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_14
cc_25 N_noxref_14_1 N_B_1 0.000991748f
cc_26 N_noxref_14_1 N_MM1_g 0.00220512f
cc_27 N_noxref_14_1 N_NET036_4 0.00163217f
cc_28 N_noxref_14_1 N_NET036_12 0.0367596f
cc_29 N_noxref_14_1 N_noxref_13_1 0.000901563f
x_PM_XOR2x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XOR2x1_ASAP7_75t_R%noxref_16
cc_30 N_noxref_16_1 N_B_1 0.00107765f
cc_31 N_noxref_16_1 N_MM5_g 0.00230453f
cc_32 N_noxref_16_1 N_NET036_4 0.00105389f
cc_33 N_noxref_16_1 N_NET019_13 0.0352749f
cc_34 N_noxref_16_1 N_noxref_14_1 0.00729301f
cc_35 N_noxref_16_1 N_noxref_15_1 0.000895648f
x_PM_XOR2x1_ASAP7_75t_R%NET019 VSS N_MM5_s N_MM4_s N_MM6_d N_MM6@2_d N_MM4@2_s
+ N_MM5@2_s N_NET019_14 N_NET019_2 N_NET019_17 N_NET019_15 N_NET019_1
+ N_NET019_3 N_NET019_13 N_NET019_16 N_NET019_4 PM_XOR2x1_ASAP7_75t_R%NET019
cc_36 N_NET019_14 N_A_21 0.000130522f
cc_37 N_NET019_14 N_A_18 0.000149977f
cc_38 N_NET019_14 N_A_17 0.000200378f
cc_39 N_NET019_14 N_A_3 0.000231432f
cc_40 N_NET019_14 N_A_16 0.000258571f
cc_41 N_NET019_14 N_A_14 0.000266269f
cc_42 N_NET019_2 N_A_2 0.000288757f
cc_43 N_NET019_17 N_A_16 0.000362002f
cc_44 N_NET019_17 N_A_18 0.000395631f
cc_45 N_NET019_15 N_MM4@2_g 0.0333616f
cc_46 N_NET019_17 N_A_22 0.000528191f
cc_47 N_NET019_1 N_A_15 0.00164041f
cc_48 N_NET019_14 N_A_2 0.000795476f
cc_49 N_NET019_15 N_A_3 0.00080383f
cc_50 N_NET019_2 N_MM4_g 0.00105734f
cc_51 N_NET019_17 N_A_24 0.00106839f
cc_52 N_NET019_3 N_MM4@2_g 0.00117005f
cc_53 N_NET019_3 N_A_18 0.00180385f
cc_54 N_NET019_17 N_A_15 0.00229606f
cc_55 N_NET019_17 N_A_25 0.00798308f
cc_56 N_NET019_14 N_MM4_g 0.0339345f
cc_57 N_NET019_13 N_MM5@2_g 6.76016e-20
cc_58 N_NET019_13 N_B_12 0.000240622f
cc_59 N_NET019_13 N_B_2 0.000367844f
cc_60 N_NET019_13 N_B_9 0.000457449f
cc_61 N_NET019_16 N_MM5@2_g 0.0335302f
cc_62 N_NET019_17 N_B_9 0.000505895f
cc_63 N_NET019_16 N_B_2 0.000770788f
cc_64 N_NET019_4 N_MM5@2_g 0.00118037f
cc_65 N_NET019_1 N_MM5_g 0.00150078f
cc_66 N_NET019_13 N_B_1 0.00208962f
cc_67 N_NET019_13 N_MM5_g 0.0341748f
cc_68 N_NET019_15 N_MM6_g 0.000435439f
cc_69 N_NET019_13 N_NET036_4 0.000594952f
cc_70 N_NET019_3 N_MM6@2_g 0.000679654f
cc_71 N_NET019_2 N_MM6_g 0.000945062f
cc_72 N_NET019_14 N_NET036_1 0.00141683f
cc_73 N_NET019_14 N_MM6_g 0.0330372f
cc_74 N_NET019_15 N_MM6@2_g 0.0348797f
x_PM_XOR2x1_ASAP7_75t_R%Y VSS Y N_MM10@2_s N_MM9_s N_MM9@2_s N_MM10_s N_MM6_s
+ N_MM6@2_s N_Y_18 N_Y_19 N_Y_4 N_Y_16 N_Y_14 N_Y_13 N_Y_1 N_Y_20 N_Y_15 N_Y_17
+ N_Y_2 N_Y_3 PM_XOR2x1_ASAP7_75t_R%Y
cc_75 N_Y_18 N_A_23 8.81211e-20
cc_76 N_Y_18 N_MM4@2_g 8.83686e-20
cc_77 N_Y_18 N_A_2 0.000207606f
cc_78 N_Y_18 N_MM4_g 9.56668e-20
cc_79 N_Y_18 N_A_17 0.000316031f
cc_80 N_Y_19 N_A_18 0.000189902f
cc_81 N_Y_4 N_MM4@2_g 0.000195563f
cc_82 N_Y_16 N_A_3 0.000218256f
cc_83 N_Y_14 N_MM4@2_g 0.00031076f
cc_84 N_Y_13 N_MM4_g 0.000324184f
cc_85 N_Y_1 N_MM4_g 0.000327264f
cc_86 N_Y_18 N_A_3 0.000360468f
cc_87 N_Y_20 N_A_18 0.000670172f
cc_88 N_Y_20 N_A_25 0.00194545f
cc_89 N_Y_18 N_A_18 0.0040947f
cc_90 N_Y_13 N_B_12 0.000119607f
cc_91 N_Y_13 N_B_9 0.00025835f
cc_92 N_Y_13 N_B_11 0.000293973f
cc_93 N_Y_13 N_B_2 0.000341826f
cc_94 N_Y_15 N_MM5@2_g 0.0342963f
cc_95 N_Y_4 N_B_9 0.000789436f
cc_96 N_Y_15 N_B_2 0.000842104f
cc_97 N_Y_18 N_B_12 0.00127557f
cc_98 N_Y_1 N_MM5_g 0.00179049f
cc_99 N_Y_4 N_MM5@2_g 0.00196314f
cc_100 N_Y_13 N_B_1 0.00234726f
cc_101 N_Y_17 N_B_12 0.00430382f
cc_102 N_Y_19 N_B_11 0.00675353f
cc_103 N_Y_13 N_MM5_g 0.034886f
cc_104 N_Y_20 N_NET036_17 0.000541528f
cc_105 N_Y_2 N_NET036_1 0.000600334f
cc_106 N_Y_16 N_MM6_g 0.03051f
cc_107 N_Y_1 N_NET036_16 0.00112373f
cc_108 N_Y_17 N_NET036_20 0.00152181f
cc_109 N_Y_3 N_MM6_g 0.00171618f
cc_110 N_Y_2 N_MM6_g 0.00212832f
cc_111 N_Y_18 N_NET036_17 0.00414889f
cc_112 N_Y_16 N_NET036_1 0.00506195f
cc_113 N_Y_17 N_NET036_16 0.0119653f
cc_114 N_Y_14 N_MM6@2_g 0.036726f
cc_115 N_Y_14 N_MM6_g 0.0685263f
cc_116 N_Y_18 N_NET019_3 0.000288099f
cc_117 N_Y_16 N_NET019_14 0.00168882f
cc_118 N_Y_16 N_NET019_15 0.000562728f
cc_119 N_Y_3 N_NET019_17 0.000686376f
cc_120 N_Y_3 N_NET019_3 0.00163213f
cc_121 N_Y_20 N_NET019_17 0.00376066f
cc_122 N_Y_3 N_NET019_2 0.00594664f
x_PM_XOR2x1_ASAP7_75t_R%NET036 VSS N_MM6_g N_MM6@2_g N_MM2_s N_MM0_s N_MM1_s
+ N_NET036_11 N_NET036_15 N_NET036_1 N_NET036_4 N_NET036_17 N_NET036_13
+ N_NET036_3 N_NET036_16 N_NET036_12 N_NET036_19 N_NET036_20
+ PM_XOR2x1_ASAP7_75t_R%NET036
cc_123 N_NET036_11 N_A_3 0.000134467f
cc_124 N_NET036_11 N_A_1 0.00107704f
cc_125 N_NET036_11 N_A_12 0.000200342f
cc_126 N_NET036_11 N_A_16 0.000216423f
cc_127 N_NET036_15 N_A_14 0.000350978f
cc_128 N_NET036_1 N_A_17 0.000361095f
cc_129 N_NET036_4 N_A_21 0.000374307f
cc_130 N_NET036_1 N_A_3 0.000375819f
cc_131 N_NET036_15 N_A_15 0.000517096f
cc_132 N_NET036_17 N_A_25 0.000553477f
cc_133 N_NET036_1 N_A_2 0.00209108f
cc_134 N_NET036_13 N_A_10 0.000711692f
cc_135 N_NET036_3 N_MM0_g 0.000976626f
cc_136 N_NET036_16 N_A_23 0.00216164f
cc_137 N_NET036_17 N_A_17 0.00253321f
cc_138 N_NET036_15 N_A_21 0.00301709f
cc_139 N_MM6@2_g N_MM4@2_g 0.00336438f
cc_140 N_MM6_g N_MM4_g 0.00341604f
cc_141 N_NET036_4 N_A_13 0.00386859f
cc_142 N_NET036_11 N_MM0_g 0.0356241f
cc_143 N_NET036_11 N_MM5_g 0.000151625f
cc_144 N_NET036_11 N_B_10 0.000784371f
cc_145 N_NET036_11 N_B_12 0.000281972f
cc_146 N_NET036_13 N_B_8 0.000449921f
cc_147 N_NET036_12 N_MM1_g 0.0161018f
cc_148 N_NET036_4 N_B_1 0.00572061f
cc_149 N_NET036_17 N_B_12 0.00065612f
cc_150 N_NET036_19 N_B_10 0.000750737f
cc_151 N_NET036_3 N_B_1 0.000834757f
cc_152 N_NET036_3 N_MM1_g 0.00144526f
cc_153 N_NET036_4 N_MM1_g 0.00289879f
cc_154 N_NET036_13 N_B_10 0.00481722f
cc_155 N_NET036_15 N_B_8 0.00580697f
cc_156 N_NET036_16 N_B_12 0.00758542f
cc_157 N_NET036_11 N_MM1_g 0.0544222f
x_PM_XOR2x1_ASAP7_75t_R%B VSS B N_MM1_g N_MM5_g N_MM5@2_g N_B_9 N_B_1 N_B_8
+ N_B_10 N_B_11 N_B_2 N_B_12 PM_XOR2x1_ASAP7_75t_R%B
cc_158 N_B_9 N_MM0_g 7.3618e-20
cc_159 N_B_1 N_MM0_g 0.00010486f
cc_160 N_B_8 N_MM0_g 0.000113357f
cc_161 N_B_9 N_A_18 0.00319957f
cc_162 N_B_1 N_A_2 0.000653227f
cc_163 N_B_8 N_A_11 0.000242425f
cc_164 N_B_1 N_A_1 0.0014196f
cc_165 N_B_1 N_A_16 0.000357919f
cc_166 N_B_10 N_A_12 0.000370564f
cc_167 N_B_1 N_A_17 0.000396773f
cc_168 N_B_11 N_A_18 0.000423919f
cc_169 N_B_1 N_A_23 0.00044829f
cc_170 N_B_10 N_A_10 0.000471084f
cc_171 N_B_1 N_A_15 0.000493497f
cc_172 N_B_8 N_A_13 0.000615838f
cc_173 N_B_2 N_A_3 0.00224312f
cc_174 N_B_8 N_A_12 0.00175969f
cc_175 N_B_12 N_A_25 0.00217005f
cc_176 N_B_1 N_A_21 0.00225076f
cc_177 N_B_12 N_A_17 0.00403854f
cc_178 N_MM5_g N_MM4_g 0.00492342f
cc_179 N_MM5@2_g N_MM4@2_g 0.00498308f
cc_180 N_MM1_g N_MM0_g 0.00527778f
x_PM_XOR2x1_ASAP7_75t_R%A VSS A N_MM0_g N_MM4_g N_MM4@2_g N_A_18 N_A_2 N_A_11
+ N_A_1 N_A_16 N_A_12 N_A_17 N_A_23 N_A_10 N_A_15 N_A_13 N_A_3 N_A_25 N_A_21
+ N_A_14 N_A_22 N_A_24 PM_XOR2x1_ASAP7_75t_R%A
*END of XOR2x1_ASAP7_75t_R.pxi
.ENDS
** Design:	XOR2x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XOR2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XOR2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XOR2x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00612301f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00470703f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%NET059 VSS 2 3 1
c1 1 VSS 0.00103195f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%NET060 VSS 2 3 1
c1 1 VSS 0.00094733f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0422838f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0049503f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00452996f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00485234f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.0310724f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0422969f
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%NET045 VSS 9 39 42 43 15 3 4 14 1 13 12 11 10 17
+ 16
c1 1 VSS 0.00186772f
c2 3 VSS 0.00615207f
c3 4 VSS 0.00751859f
c4 9 VSS 0.0422073f
c5 10 VSS 0.00475297f
c6 11 VSS 0.00592487f
c7 12 VSS 0.00169687f
c8 13 VSS 0.00547947f
c9 14 VSS 0.00187733f
c10 15 VSS 0.00171904f
c11 16 VSS 0.000464214f
c12 17 VSS 0.000492684f
r1 43 41 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r2 37 41 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2160 $X2=0.3925 $Y2=0.2160
r3 11 37 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2160 $X2=0.3780 $Y2=0.2160
r4 42 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2160 $X2=0.3635 $Y2=0.2160
r5 39 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r6 10 38 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.0675 $X2=0.3385 $Y2=0.0675
r7 4 37 17.0927 $w=2.02e-08 $l=2.9e-08 $layer=LISD $thickness=2.7e-08 $X=0.3780
+ $Y=0.1870 $X2=0.3780 $Y2=0.2160
r8 3 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3115 $Y=0.0675
+ $X2=0.3110 $Y2=0.0930
r9 33 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3745 $Y=0.1980
+ $X2=0.3780 $Y2=0.2160
r10 32 33 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.1980 $X2=0.3745 $Y2=0.1980
r11 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.3645 $Y2=0.1980
r12 15 17 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.1980 $X2=0.3110 $Y2=0.1980
r13 15 31 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r14 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.0930 $X2=0.3110 $Y2=0.1245
r15 26 28 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.1565 $X2=0.3110 $Y2=0.1245
r16 14 17 3.94987 $w=1.50455e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3110 $Y=0.1760 $X2=0.3110 $Y2=0.1980
r17 14 26 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.1760 $X2=0.3110 $Y2=0.1565
r18 17 25 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3110 $Y=0.1980 $X2=0.2905 $Y2=0.1980
r19 24 25 18.422 $w=1.3e-08 $l=7.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2115
+ $Y=0.1980 $X2=0.2905 $Y2=0.1980
r20 23 24 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.2115 $Y2=0.1980
r21 22 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1125
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r22 13 16 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.1980 $X2=0.0810 $Y2=0.1980
r23 13 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1125 $Y2=0.1980
r24 16 21 4.9968 $w=1.60947e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.1980 $X2=0.0810 $Y2=0.1695
r25 20 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1470 $X2=0.0810 $Y2=0.1695
r26 19 20 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1470
r27 12 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r28 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r29 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r30 3 10 1e-05
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%Y VSS 21 16 17 28 29 9 7 8 10 11 2 1
c1 1 VSS 0.0104224f
c2 2 VSS 0.00998413f
c3 7 VSS 0.00447474f
c4 8 VSS 0.00448715f
c5 9 VSS 0.00842429f
c6 10 VSS 0.00876967f
c7 11 VSS 0.00702289f
c8 12 VSS 0.00344628f
c9 13 VSS 0.00336385f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r6 10 13 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5265 $Y=0.2340 $X2=0.5670 $Y2=0.2340
r7 10 25 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r8 13 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.2340 $X2=0.5670 $Y2=0.2160
r9 22 23 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1775 $X2=0.5670 $Y2=0.2160
r10 21 22 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1475 $X2=0.5670 $Y2=0.1775
r11 21 20 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1475 $X2=0.5670 $Y2=0.1330
r12 11 12 9.07762 $w=1.49174e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0820 $X2=0.5670 $Y2=0.0360
r13 11 20 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0820 $X2=0.5670 $Y2=0.1330
r14 12 19 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5265 $Y2=0.0360
r15 9 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5265 $Y2=0.0360
r16 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r17 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r18 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r19 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r20 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%NET049 VSS 12 13 19 7 8 1 9 2
c1 1 VSS 0.00722435f
c2 2 VSS 0.0075559f
c3 7 VSS 0.00340297f
c4 8 VSS 0.00371023f
c5 9 VSS 0.0132415f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r2 19 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r3 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0360
r4 15 16 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1665
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r5 14 15 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1665 $Y2=0.0360
r6 9 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r7 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r8 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r9 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r10 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r11 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%A VSS 23 3 4 5 1 6
c1 1 VSS 0.00930203f
c2 3 VSS 0.0465406f
c3 4 VSS 0.0358075f
c4 5 VSS 0.00378204f
c5 6 VSS 0.0038495f
r1 6 22 3.3086 $w=1.53377e-08 $l=1.92e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3510 $Y2=0.0912
r2 3 17 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 23 24 2.85657 $w=1.3e-08 $l=1.22e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1020 $X2=0.3510 $Y2=0.1142
r4 23 22 2.50679 $w=1.3e-08 $l=1.08e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1020 $X2=0.3510 $Y2=0.0912
r5 5 20 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1265 $X2=0.3510 $Y2=0.1350
r6 5 24 2.85657 $w=1.3e-08 $l=1.23e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1265 $X2=0.3510 $Y2=0.1142
r7 15 17 10.5547 $w=1.466e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r8 14 15 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2015 $Y2=0.1350
r9 13 14 96.7394 $w=9.3e-09 $l=4.15e-08 $layer=LIG $thickness=4.8e-08 $X=0.2575
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r10 12 13 97.9049 $w=9.3e-09 $l=4.2e-08 $layer=LIG $thickness=4.8e-08 $X=0.2995
+ $Y=0.1350 $X2=0.2575 $Y2=0.1350
r11 11 12 57.1112 $w=9.3e-09 $l=2.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.2995 $Y2=0.1350
r12 10 11 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r13 9 19 1.40189 $w=1.265e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3605
+ $Y=0.1350 $X2=0.3615 $Y2=0.1350
r14 8 9 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3605 $Y2=0.1350
r15 8 20 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r16 1 8 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r17 1 10 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3415 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r18 4 8 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r19 4 10 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r20 4 19 1.4802 $w=2.16633e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3615 $Y2=0.1350
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%B VSS 24 5 6 14 2 9 15 8 1 7 10 11 12 17 16
c1 1 VSS 0.0054021f
c2 2 VSS 0.00591124f
c3 5 VSS 0.0824518f
c4 6 VSS 0.0826255f
c5 7 VSS 0.00193943f
c6 8 VSS 0.00322441f
c7 9 VSS 0.00122904f
c8 10 VSS 0.0141464f
c9 11 VSS 0.00359118f
c10 12 VSS 0.00127876f
c11 13 VSS 0.00294406f
c12 14 VSS 0.0010295f
c13 15 VSS 0.00116737f
c14 16 VSS 0.00337212f
c15 17 VSS 0.00155272f
r1 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r2 5 1 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 38 39 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1235 $X2=0.1350 $Y2=0.1350
r4 7 12 4.41382 $w=1.63923e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1040 $X2=0.1350 $Y2=0.0780
r5 7 38 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1040 $X2=0.1350 $Y2=0.1235
r6 12 37 10.4768 $w=1.38654e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0780 $X2=0.1870 $Y2=0.0780
r7 8 14 3.92057 $w=1.38108e-08 $l=2.5224e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2455 $Y=0.0780 $X2=0.2700 $Y2=0.0720
r8 8 37 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2455
+ $Y=0.0780 $X2=0.1870 $Y2=0.0780
r9 14 35 1.0057 $w=1.55e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0720 $X2=0.2700 $Y2=0.0660
r10 9 13 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0360
r11 9 35 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0540 $X2=0.2700 $Y2=0.0660
r12 13 34 3.13128 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.0360 $X2=0.2905 $Y2=0.0360
r13 33 34 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.0360 $X2=0.2905 $Y2=0.0360
r14 32 33 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.0360 $X2=0.3110 $Y2=0.0360
r15 31 32 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3610
+ $Y=0.0360 $X2=0.3310 $Y2=0.0360
r16 30 31 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3855
+ $Y=0.0360 $X2=0.3610 $Y2=0.0360
r17 10 16 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4065 $Y=0.0360 $X2=0.4310 $Y2=0.0360
r18 10 30 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4065
+ $Y=0.0360 $X2=0.3855 $Y2=0.0360
r19 16 29 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.0360 $X2=0.4310 $Y2=0.0540
r20 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.0720 $X2=0.4310 $Y2=0.0540
r21 27 28 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1000 $X2=0.4310 $Y2=0.0720
r22 11 17 1.24985 $w=1.57419e-08 $l=7.7e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4310 $Y=0.1225 $X2=0.4310 $Y2=0.1302
r23 11 27 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1225 $X2=0.4310 $Y2=0.1000
r24 24 17 0.484711 $w=1.8e-08 $l=4.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1350 $X2=0.4310 $Y2=0.1302
r25 24 23 0.983781 $w=1.35556e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4310 $Y=0.1350 $X2=0.4180 $Y2=0.1350
r26 22 23 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4180 $Y2=0.1350
r27 21 22 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r28 15 21 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1350 $X2=0.3940 $Y2=0.1350
r29 6 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r30 2 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_XOR2x2_ASAP7_75t_R%XOR VSS 12 13 50 55 59 4 19 18 5 15 24 3 14 17 16
+ 1 22 20 21 26 25
c1 1 VSS 0.00708864f
c2 3 VSS 0.00573441f
c3 4 VSS 0.00813559f
c4 5 VSS 0.00574941f
c5 12 VSS 0.0803064f
c6 13 VSS 0.0808523f
c7 14 VSS 0.00458849f
c8 15 VSS 0.00582924f
c9 16 VSS 0.00502874f
c10 17 VSS 0.00753845f
c11 18 VSS 0.0365668f
c12 19 VSS 0.000693528f
c13 20 VSS 0.00116471f
c14 21 VSS 0.00201757f
c15 22 VSS 0.0065816f
c16 23 VSS 0.00341479f
c17 24 VSS 0.000742528f
c18 25 VSS 0.00299698f
c19 26 VSS 0.000442752f
r1 59 58 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r2 14 58 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r3 3 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r4 56 57 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r5 22 53 3.71668 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0570
r6 22 56 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r7 55 54 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r8 15 54 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r9 52 53 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0950 $X2=0.0270 $Y2=0.0570
r10 51 52 16.0901 $w=1.3e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1640 $X2=0.0270 $Y2=0.0950
r11 17 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2160 $X2=0.0270 $Y2=0.2340
r12 17 51 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2160 $X2=0.0270 $Y2=0.1640
r13 16 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r14 50 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r15 4 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r16 23 45 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r17 5 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2160
+ $X2=0.2160 $Y2=0.2340
r18 45 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r19 44 46 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r20 42 43 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r21 41 42 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1395
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r22 41 44 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1395
+ $Y=0.2340 $X2=0.0675 $Y2=0.2340
r23 40 43 22.9692 $w=1.3e-08 $l=9.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4070
+ $Y=0.2340 $X2=0.3085 $Y2=0.2340
r24 18 25 0.56619 $w=1.77368e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4225 $Y=0.2340 $X2=0.4320 $Y2=0.2340
r25 18 40 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4225
+ $Y=0.2340 $X2=0.4070 $Y2=0.2340
r26 19 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2160 $X2=0.4320 $Y2=0.1980
r27 19 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2160 $X2=0.4320 $Y2=0.2340
r28 24 39 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.1980 $X2=0.4565 $Y2=0.1980
r29 20 26 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4745 $Y=0.1980 $X2=0.4860 $Y2=0.1980
r30 20 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4745
+ $Y=0.1980 $X2=0.4565 $Y2=0.1980
r31 26 37 3.48106 $w=1.70091e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.1980 $X2=0.4860 $Y2=0.1760
r32 13 33 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r33 36 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1535 $X2=0.4860 $Y2=0.1760
r34 35 36 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1350 $X2=0.4860 $Y2=0.1535
r35 21 35 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1225 $X2=0.4860 $Y2=0.1350
r36 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r37 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r38 30 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4860 $Y=0.1350
+ $X2=0.4860 $Y2=0.1350
r39 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r40 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r41 1 28 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4485 $Y2=0.1350
r42 1 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r43 12 28 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4590 $Y=0.1350 $X2=0.4485 $Y2=0.1350
r44 12 29 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r45 3 14 1e-05
r46 4 15 1e-05
.ends


*
.SUBCKT XOR2x2_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM0_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 VSS N_MM12_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13@2 VSS N_MM12@2_g N_MM13@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM5_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM4_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM12 VDD N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12@2 VDD N_MM12@2_g N_MM12@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XOR2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XOR2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XOR2x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_13
cc_1 N_noxref_13_1 N_NET045_3 0.00100712f
cc_2 N_noxref_13_1 N_A_1 0.00108511f
cc_3 N_noxref_13_1 N_MM4_g 0.00229947f
cc_4 N_noxref_13_1 N_NET049_8 0.0352251f
x_PM_XOR2x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_15
cc_5 N_noxref_15_1 N_NET045_3 0.00158325f
cc_6 N_noxref_15_1 N_NET045_10 0.0366845f
cc_7 N_noxref_15_1 N_A_1 0.00100321f
cc_8 N_noxref_15_1 N_MM0_g 0.00228811f
cc_9 N_noxref_15_1 N_noxref_13_1 0.00730784f
x_PM_XOR2x2_ASAP7_75t_R%NET059 VSS N_MM11_d N_MM10_s N_NET059_1
+ PM_XOR2x2_ASAP7_75t_R%NET059
cc_10 N_NET059_1 N_MM5_g 0.0173114f
cc_11 N_NET059_1 N_MM4_g 0.0173033f
x_PM_XOR2x2_ASAP7_75t_R%NET060 VSS N_MM2_s N_MM3_d N_NET060_1
+ PM_XOR2x2_ASAP7_75t_R%NET060
cc_12 N_NET060_1 N_MM1_g 0.0172999f
cc_13 N_NET060_1 N_MM0_g 0.0174599f
x_PM_XOR2x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_17
cc_14 N_noxref_17_1 N_MM12@2_g 0.00147155f
cc_15 N_noxref_17_1 N_Y_7 0.000835897f
x_PM_XOR2x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_14
cc_16 N_noxref_14_1 N_A_1 0.00114473f
cc_17 N_noxref_14_1 N_MM4_g 0.00235882f
cc_18 N_noxref_14_1 N_XOR_16 0.0370192f
cc_19 N_noxref_14_1 N_noxref_13_1 0.000896035f
x_PM_XOR2x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_12
cc_20 N_noxref_12_1 N_MM6_g 0.0014537f
cc_21 N_noxref_12_1 N_XOR_17 0.000325763f
cc_22 N_noxref_12_1 N_XOR_4 0.000508146f
cc_23 N_noxref_12_1 N_XOR_15 0.0377831f
cc_24 N_noxref_12_1 N_noxref_11_1 0.00176442f
x_PM_XOR2x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_11
cc_25 N_noxref_11_1 N_MM6_g 0.00145195f
cc_26 N_noxref_11_1 N_XOR_17 0.000326924f
cc_27 N_noxref_11_1 N_XOR_3 0.000509729f
cc_28 N_noxref_11_1 N_XOR_14 0.0375217f
x_PM_XOR2x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_16
cc_29 N_noxref_16_1 N_NET045_11 0.00048983f
cc_30 N_noxref_16_1 N_A_1 0.00141509f
cc_31 N_noxref_16_1 N_MM0_g 0.0043005f
cc_32 N_noxref_16_1 N_XOR_16 0.000553163f
cc_33 N_noxref_16_1 N_noxref_14_1 0.00751029f
cc_34 N_noxref_16_1 N_noxref_15_1 0.000968181f
x_PM_XOR2x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_XOR2x2_ASAP7_75t_R%noxref_18
cc_35 N_noxref_18_1 N_MM12@2_g 0.00147742f
cc_36 N_noxref_18_1 N_Y_8 0.000829038f
cc_37 N_noxref_18_1 N_noxref_17_1 0.00176783f
x_PM_XOR2x2_ASAP7_75t_R%NET045 VSS N_MM6_g N_MM2_d N_MM0_d N_MM1_d N_NET045_15
+ N_NET045_3 N_NET045_4 N_NET045_14 N_NET045_1 N_NET045_13 N_NET045_12
+ N_NET045_11 N_NET045_10 N_NET045_17 N_NET045_16 PM_XOR2x2_ASAP7_75t_R%NET045
x_PM_XOR2x2_ASAP7_75t_R%Y VSS Y N_MM13_s N_MM13@2_s N_MM12_s N_MM12@2_s N_Y_9
+ N_Y_7 N_Y_8 N_Y_10 N_Y_11 N_Y_2 N_Y_1 PM_XOR2x2_ASAP7_75t_R%Y
cc_38 N_Y_9 N_B_11 0.00089391f
cc_39 N_Y_9 N_B_16 0.00252019f
cc_40 N_Y_7 N_XOR_21 0.000295021f
cc_41 N_Y_7 N_XOR_26 0.0003675f
cc_42 N_Y_7 N_XOR_25 0.000384209f
cc_43 N_Y_7 N_XOR_1 0.00075581f
cc_44 N_Y_8 N_MM12_g 0.0308086f
cc_45 N_Y_10 N_XOR_20 0.000968341f
cc_46 N_Y_11 N_XOR_1 0.00129167f
cc_47 N_Y_2 N_XOR_21 0.00173853f
cc_48 N_Y_1 N_MM12_g 0.00197203f
cc_49 N_Y_2 N_MM12_g 0.00259315f
cc_50 N_Y_10 N_XOR_26 0.00315499f
cc_51 N_Y_8 N_XOR_1 0.00424081f
cc_52 N_Y_7 N_MM12@2_g 0.0370799f
cc_53 N_Y_7 N_MM12_g 0.0682531f
x_PM_XOR2x2_ASAP7_75t_R%NET049 VSS N_MM6_s N_MM5_d N_MM4_d N_NET049_7
+ N_NET049_8 N_NET049_1 N_NET049_9 N_NET049_2 PM_XOR2x2_ASAP7_75t_R%NET049
cc_54 N_NET049_7 N_NET045_3 0.000413148f
cc_55 N_NET049_8 N_NET045_3 0.000569249f
cc_56 N_NET049_7 N_NET045_1 0.000633311f
cc_57 N_NET049_1 N_MM6_g 0.000880429f
cc_58 N_NET049_7 N_MM6_g 0.0343641f
cc_59 N_NET049_7 N_B_8 0.000405384f
cc_60 N_NET049_1 N_B_7 0.000505193f
cc_61 N_NET049_7 N_B_1 0.000738973f
cc_62 N_NET049_9 N_B_12 0.000949914f
cc_63 N_NET049_2 N_B_8 0.00106804f
cc_64 N_NET049_1 N_MM5_g 0.00124475f
cc_65 N_NET049_9 N_B_8 0.00718587f
cc_66 N_NET049_7 N_MM5_g 0.0347453f
cc_67 N_NET049_2 N_MM4_g 0.00153065f
cc_68 N_NET049_8 N_A_1 0.00218124f
cc_69 N_NET049_8 N_MM4_g 0.033957f
cc_70 N_NET049_1 N_XOR_14 0.00112737f
cc_71 N_NET049_9 N_XOR_22 0.000883403f
cc_72 N_NET049_1 N_XOR_3 0.0040476f
x_PM_XOR2x2_ASAP7_75t_R%A VSS A N_MM4_g N_MM0_g N_A_5 N_A_1 N_A_6
+ PM_XOR2x2_ASAP7_75t_R%A
cc_73 N_A_5 N_NET045_10 0.000292882f
cc_74 N_MM0_g N_NET045_4 0.000570275f
cc_75 N_A_5 N_NET045_3 0.000641839f
cc_76 N_A_1 N_NET045_13 0.000773961f
cc_77 N_A_6 N_NET045_14 0.000807758f
cc_78 N_A_1 N_NET045_14 0.000854188f
cc_79 N_A_5 N_NET045_15 0.000959159f
cc_80 N_MM0_g N_NET045_3 0.00321465f
cc_81 N_MM0_g N_NET045_11 0.0109106f
cc_82 N_A_1 N_NET045_3 0.00511404f
cc_83 N_A_5 N_NET045_14 0.00756499f
cc_84 N_MM0_g N_NET045_10 0.0498741f
cc_85 N_A_1 N_MM1_g 0.000809768f
cc_86 N_A_1 N_B_8 0.000474154f
cc_87 N_A_1 N_B_1 0.000480419f
cc_88 N_A_1 N_B_2 0.00138106f
cc_89 N_A_6 N_B_11 0.000621691f
cc_90 N_A_1 N_B_14 0.00204088f
cc_91 N_A_5 N_B_15 0.00253256f
cc_92 N_MM4_g N_MM5_g 0.00490625f
cc_93 N_A_6 N_B_10 0.00507407f
cc_94 N_MM0_g N_MM1_g 0.00748899f
x_PM_XOR2x2_ASAP7_75t_R%B VSS B N_MM5_g N_MM1_g N_B_14 N_B_2 N_B_9 N_B_15 N_B_8
+ N_B_1 N_B_7 N_B_10 N_B_11 N_B_12 N_B_17 N_B_16 PM_XOR2x2_ASAP7_75t_R%B
cc_95 N_MM1_g N_NET045_15 0.000288361f
cc_96 N_B_14 N_NET045_3 0.000358124f
cc_97 N_B_2 N_NET045_4 0.00038405f
cc_98 N_B_9 N_NET045_14 0.000448828f
cc_99 N_MM1_g N_NET045_4 0.000507798f
cc_100 N_B_15 N_NET045_15 0.000789448f
cc_101 N_B_8 N_NET045_3 0.000873352f
cc_102 N_B_1 N_NET045_1 0.00192212f
cc_103 N_B_7 N_NET045_13 0.00156726f
cc_104 N_B_10 N_NET045_3 0.00162945f
cc_105 N_B_10 N_NET045_14 0.00164087f
cc_106 N_B_7 N_NET045_12 0.00285703f
cc_107 N_B_14 N_NET045_14 0.00303243f
cc_108 N_MM5_g N_MM6_g 0.00336305f
cc_109 N_MM1_g N_NET045_11 0.0260681f
x_PM_XOR2x2_ASAP7_75t_R%XOR VSS N_MM12_g N_MM12@2_g N_MM10_d N_MM9_d N_MM6_d
+ N_XOR_4 N_XOR_19 N_XOR_18 N_XOR_5 N_XOR_15 N_XOR_24 N_XOR_3 N_XOR_14 N_XOR_17
+ N_XOR_16 N_XOR_1 N_XOR_22 N_XOR_20 N_XOR_21 N_XOR_26 N_XOR_25
+ PM_XOR2x2_ASAP7_75t_R%XOR
cc_110 N_XOR_4 N_MM6_g 0.00158853f
cc_111 N_XOR_19 N_MM6_g 0.00020738f
cc_112 N_XOR_18 N_NET045_14 0.000284539f
cc_113 N_XOR_5 N_NET045_13 0.00154128f
cc_114 N_XOR_15 N_MM6_g 0.0159003f
cc_115 N_XOR_18 N_NET045_4 0.000961865f
cc_116 N_XOR_24 N_NET045_15 0.000483699f
cc_117 N_XOR_4 N_NET045_1 0.000911857f
cc_118 N_XOR_3 N_MM6_g 0.00106956f
cc_119 N_XOR_18 N_NET045_17 0.00118309f
cc_120 N_XOR_14 N_NET045_1 0.00163646f
cc_121 N_XOR_18 N_NET045_16 0.00172118f
cc_122 N_XOR_18 N_NET045_15 0.00289156f
cc_123 N_XOR_17 N_NET045_12 0.00469106f
cc_124 N_XOR_18 N_NET045_13 0.0212429f
cc_125 N_XOR_14 N_MM6_g 0.0541978f
cc_126 N_XOR_16 N_MM1_g 9.60431e-20
cc_127 N_XOR_4 N_MM1_g 0.000110053f
cc_128 N_XOR_15 N_MM1_g 0.0001143f
cc_129 N_XOR_1 N_MM1_g 0.000195129f
cc_130 N_XOR_24 N_MM1_g 0.000202259f
cc_131 N_XOR_5 N_MM1_g 0.000208758f
cc_132 N_XOR_22 N_B_12 0.000229818f
cc_133 N_XOR_17 N_B_7 0.000269117f
cc_134 N_XOR_1 N_B_17 0.00027354f
cc_135 N_XOR_5 N_MM5_g 0.000305078f
cc_136 N_XOR_18 N_B_7 0.000328522f
cc_137 N_XOR_14 N_MM5_g 0.000342595f
cc_138 N_XOR_20 N_B_17 0.000368575f
cc_139 N_XOR_3 N_B_7 0.000368729f
cc_140 N_XOR_21 N_B_11 0.000788352f
cc_141 N_XOR_1 N_B_2 0.00110568f
cc_142 N_XOR_21 N_B_17 0.00168844f
cc_143 N_XOR_24 N_B_17 0.00203292f
cc_144 N_MM12_g N_MM1_g 0.0038854f
cc_145 N_XOR_24 N_A_5 0.000200215f
cc_146 N_XOR_5 N_MM4_g 0.00180505f
cc_147 N_XOR_16 N_A_1 0.00246501f
cc_148 N_XOR_16 N_MM4_g 0.0364995f
*END of XOR2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	XOR2xp5_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XOR2xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XOR2xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00541371f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00460471f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00624318f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00478038f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00485927f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0315616f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%Y VSS 25 18 29 33 1 10 2 3 13 12 14 11 15
c1 1 VSS 0.00661774f
c2 2 VSS 0.00791769f
c3 3 VSS 0.00595601f
c4 10 VSS 0.00366401f
c5 11 VSS 0.00355773f
c6 12 VSS 0.00245422f
c7 13 VSS 0.0177615f
c8 14 VSS 0.00313311f
c9 15 VSS 0.00547636f
c10 16 VSS 0.00281387f
r1 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r2 33 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r3 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r4 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r5 15 27 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r6 15 31 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r7 11 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r8 29 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r9 26 27 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4590 $Y2=0.2160
r10 25 26 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1060 $X2=0.4590 $Y2=0.1780
r11 14 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r12 25 14 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1060 $X2=0.4590 $Y2=0.0540
r13 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r14 16 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4455 $Y2=0.0360
r15 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r16 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r17 21 22 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3465
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r18 20 21 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3465 $Y2=0.0360
r19 13 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r20 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0540
+ $X2=0.2700 $Y2=0.0360
r21 18 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r22 10 17 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r23 1 10 1e-05
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%NET047 VSS 2 3 1
c1 1 VSS 0.00100786f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3240 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.0675 $X2=0.3240 $Y2=0.0675
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0321379f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%NET048 VSS 2 3 1
c1 1 VSS 0.00093787f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1080 $Y2=0.2025
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0419889f
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%NET019 VSS 11 18 19 8 1 2 9 7
c1 1 VSS 0.00700365f
c2 2 VSS 0.00708466f
c3 7 VSS 0.00370637f
c4 8 VSS 0.00338573f
c5 9 VSS 0.0113861f
r1 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 2 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 18 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 2 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3780 $Y2=0.2340
r6 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.2340 $X2=0.3780 $Y2=0.2340
r7 13 14 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3195
+ $Y=0.2340 $X2=0.3645 $Y2=0.2340
r8 12 13 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3195 $Y2=0.2340
r9 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r10 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r11 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r12 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r13 1 7 1e-05
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%B VSS 21 3 4 1 6 7 5
c1 1 VSS 0.00869522f
c2 3 VSS 0.0355556f
c3 4 VSS 0.0461873f
c4 5 VSS 0.00372095f
c5 6 VSS 0.00346923f
c6 7 VSS 0.00369725f
r1 6 24 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 7 23 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 19 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 22 24 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1435 $X2=0.1350 $Y2=0.1665
r5 21 22 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1435
r6 21 5 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1265
r7 5 23 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1035
r8 17 19 10.5547 $w=1.466e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 16 17 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2845 $Y2=0.1350
r10 15 16 96.7394 $w=9.3e-09 $l=4.15e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2285 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r11 14 15 97.9049 $w=9.3e-09 $l=4.2e-08 $layer=LIG $thickness=4.8e-08 $X=0.1865
+ $Y=0.1350 $X2=0.2285 $Y2=0.1350
r12 13 14 57.1112 $w=9.3e-09 $l=2.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1865 $Y2=0.1350
r13 12 13 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r14 10 12 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1445 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r15 9 10 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r16 21 9 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r17 1 9 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r18 1 11 1.40189 $w=1.265e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1245 $Y2=0.1350
r19 3 9 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r20 3 11 1.4802 $w=2.16633e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1245 $Y2=0.1350
r21 3 12 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%A VSS 25 5 6 1 12 9 2 16 10 7 13 17 18
c1 1 VSS 0.00556457f
c2 2 VSS 0.00412903f
c3 5 VSS 0.0715445f
c4 6 VSS 0.0825556f
c5 7 VSS 0.0110363f
c6 8 VSS 0.00737687f
c7 9 VSS 0.00204822f
c8 10 VSS 0.0186816f
c9 11 VSS 0.000355211f
c10 12 VSS 0.00415084f
c11 13 VSS 0.00347077f
c12 14 VSS 0.00186784f
c13 15 VSS 0.00472596f
c14 16 VSS 0.000415132f
c15 17 VSS 0.0029344f
c16 18 VSS 0.000832674f
r1 2 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r2 6 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 41 42 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1465
r4 13 18 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1690 $X2=0.3510 $Y2=0.1980
r5 13 42 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1690 $X2=0.3510 $Y2=0.1465
r6 18 39 10.4768 $w=1.38654e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.2990 $Y2=0.1980
r7 12 16 4.22671 $w=1.43953e-08 $l=2.4683e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2405 $Y=0.1980 $X2=0.2160 $Y2=0.2010
r8 12 39 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2405
+ $Y=0.1980 $X2=0.2990 $Y2=0.1980
r9 11 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2160 $X2=0.2160 $Y2=0.2340
r10 11 16 2.71097 $w=1.5e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2160 $X2=0.2160 $Y2=0.2010
r11 17 37 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.2340 $X2=0.1935 $Y2=0.2340
r12 36 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.2340 $X2=0.1935 $Y2=0.2340
r13 35 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1710 $Y2=0.2340
r14 34 35 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1250
+ $Y=0.2340 $X2=0.1530 $Y2=0.2340
r15 33 34 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1000
+ $Y=0.2340 $X2=0.1250 $Y2=0.2340
r16 32 33 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0860
+ $Y=0.2340 $X2=0.1000 $Y2=0.2340
r17 10 15 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.2340 $X2=0.0270 $Y2=0.2340
r18 10 32 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.2340 $X2=0.0860 $Y2=0.2340
r19 15 31 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.2340 $X2=0.0270 $Y2=0.2160
r20 30 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1980 $X2=0.0270 $Y2=0.2160
r21 8 14 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r22 8 30 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1665 $X2=0.0270 $Y2=0.1980
r23 7 14 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r24 25 9 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r25 9 14 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r26 25 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r27 21 23 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r28 1 20 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r29 1 21 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r30 5 20 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r31 5 21 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_XOR2xp5_ASAP7_75t_R%NET036 VSS 9 38 41 42 14 10 4 3 12 1 15 16 11 13
+ 18 19
c1 1 VSS 0.00167816f
c2 3 VSS 0.00889377f
c3 4 VSS 0.00619883f
c4 9 VSS 0.0421499f
c5 10 VSS 0.00581069f
c6 11 VSS 0.0046823f
c7 12 VSS 0.0072376f
c8 13 VSS 0.000786085f
c9 14 VSS 0.0019145f
c10 15 VSS 0.00681309f
c11 16 VSS 0.00157342f
c12 17 VSS 0.00274831f
c13 18 VSS 0.000512152f
c14 19 VSS 0.000425872f
r1 42 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r2 3 40 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0540 $X2=0.1225 $Y2=0.0540
r3 10 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0540 $X2=0.1080 $Y2=0.0540
r4 41 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0540 $X2=0.0935 $Y2=0.0540
r5 3 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0540
+ $X2=0.1120 $Y2=0.0360
r6 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.2025 $X2=0.1600 $Y2=0.2025
r7 38 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1475 $Y2=0.2025
r8 32 33 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r9 12 17 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1710 $Y2=0.0360
r10 12 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1305 $Y2=0.0360
r11 4 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1745 $Y=0.2025
+ $X2=0.1710 $Y2=0.1800
r12 29 30 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1455 $X2=0.1710 $Y2=0.1800
r13 14 18 5.4656 $w=1.45789e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.1005 $X2=0.1710 $Y2=0.0720
r14 14 29 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1005 $X2=0.1710 $Y2=0.1455
r15 13 18 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0540 $X2=0.1710 $Y2=0.0720
r16 13 17 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0540 $X2=0.1710 $Y2=0.0360
r17 18 28 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0720 $X2=0.1935 $Y2=0.0720
r18 27 28 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.0720 $X2=0.1935 $Y2=0.0720
r19 26 27 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2990
+ $Y=0.0720 $X2=0.2315 $Y2=0.0720
r20 25 26 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.2990 $Y2=0.0720
r21 24 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3735
+ $Y=0.0720 $X2=0.3510 $Y2=0.0720
r22 15 19 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3915 $Y=0.0720 $X2=0.4050 $Y2=0.0720
r23 15 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.0720 $X2=0.3735 $Y2=0.0720
r24 19 23 4.9968 $w=1.60947e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.0720 $X2=0.4050 $Y2=0.1005
r25 16 21 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1230 $X2=0.4050 $Y2=0.1350
r26 16 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1230 $X2=0.4050 $Y2=0.1005
r27 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r28 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends


*
.SUBCKT XOR2xp5_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM0 VSS N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 VSS N_MM1_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM10_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VSS N_MM11_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 VSS N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM0_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM1_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 VDD N_MM10_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 VDD N_MM11_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM9_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XOR2xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XOR2xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XOR2xp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_B_1 0.00113715f
cc_2 N_noxref_14_1 N_MM10_g 0.0023561f
cc_3 N_noxref_14_1 N_Y_10 0.0365466f
cc_4 N_noxref_14_1 N_noxref_12_1 0.00749033f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_13
cc_5 N_noxref_13_1 N_B_1 0.000991179f
cc_6 N_noxref_13_1 N_MM1_g 0.00228133f
cc_7 N_noxref_13_1 N_NET036_4 0.00158701f
cc_8 N_noxref_13_1 N_NET036_11 0.0368277f
cc_9 N_noxref_13_1 N_noxref_12_1 0.000965398f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_15
cc_10 N_noxref_15_1 N_B_1 0.00108047f
cc_11 N_noxref_15_1 N_MM10_g 0.00230394f
cc_12 N_noxref_15_1 N_NET036_4 0.00100694f
cc_13 N_noxref_15_1 N_NET019_7 0.035109f
cc_14 N_noxref_15_1 N_noxref_13_1 0.00731502f
cc_15 N_noxref_15_1 N_noxref_14_1 0.000895268f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_16
cc_16 N_noxref_16_1 N_MM9_g 0.00145722f
cc_17 N_noxref_16_1 N_Y_11 0.0384714f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_17
cc_18 N_noxref_17_1 N_MM9_g 0.00145624f
cc_19 N_noxref_17_1 N_Y_12 0.0383331f
cc_20 N_noxref_17_1 N_noxref_16_1 0.00177384f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_12
cc_21 N_noxref_12_1 N_B_1 0.00138916f
cc_22 N_noxref_12_1 N_MM1_g 0.00431442f
cc_23 N_noxref_12_1 N_NET036_10 0.000512876f
x_PM_XOR2xp5_ASAP7_75t_R%Y VSS Y N_MM10_s N_MM9_s N_MM6_s N_Y_1 N_Y_10 N_Y_2
+ N_Y_3 N_Y_13 N_Y_12 N_Y_14 N_Y_11 N_Y_15 PM_XOR2xp5_ASAP7_75t_R%Y
cc_24 N_Y_1 N_MM10_g 0.00181305f
cc_25 N_Y_10 N_B_1 0.00237744f
cc_26 N_Y_10 N_MM10_g 0.035978f
cc_27 N_Y_2 N_NET036_1 0.000851689f
cc_28 N_Y_3 N_MM9_g 0.00107046f
cc_29 N_Y_1 N_NET036_15 0.00121723f
cc_30 N_Y_2 N_MM9_g 0.0014052f
cc_31 N_Y_13 N_NET036_19 0.00145324f
cc_32 N_Y_12 N_NET036_1 0.00157841f
cc_33 N_Y_14 N_NET036_16 0.00447797f
cc_34 N_Y_12 N_MM9_g 0.0152006f
cc_35 N_Y_13 N_NET036_15 0.0136871f
cc_36 N_Y_11 N_MM9_g 0.0553589f
cc_37 N_Y_15 N_NET019_9 0.000746918f
cc_38 N_Y_3 N_NET019_2 0.00516339f
x_PM_XOR2xp5_ASAP7_75t_R%NET047 VSS N_MM10_d N_MM11_s N_NET047_1
+ PM_XOR2xp5_ASAP7_75t_R%NET047
cc_39 N_NET047_1 N_MM11_g 0.0172237f
cc_40 N_NET047_1 N_MM10_g 0.0174148f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_10
cc_41 N_noxref_10_1 N_MM0_g 0.00466932f
x_PM_XOR2xp5_ASAP7_75t_R%NET048 VSS N_MM3_s N_MM2_d N_NET048_1
+ PM_XOR2xp5_ASAP7_75t_R%NET048
cc_42 N_NET048_1 N_MM0_g 0.0174958f
cc_43 N_NET048_1 N_MM1_g 0.0174003f
x_PM_XOR2xp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XOR2xp5_ASAP7_75t_R%noxref_11
cc_44 N_noxref_11_1 N_MM0_g 0.00263963f
cc_45 N_noxref_11_1 N_noxref_10_1 0.00185044f
x_PM_XOR2xp5_ASAP7_75t_R%NET019 VSS N_MM5_s N_MM4_s N_MM6_d N_NET019_8
+ N_NET019_1 N_NET019_2 N_NET019_9 N_NET019_7 PM_XOR2xp5_ASAP7_75t_R%NET019
cc_46 N_NET019_8 N_A_17 0.000475495f
cc_47 N_NET019_1 N_A_12 0.00156078f
cc_48 N_NET019_2 N_A_13 0.000600592f
cc_49 N_NET019_8 N_A_2 0.000778754f
cc_50 N_NET019_2 N_MM11_g 0.00129278f
cc_51 N_NET019_9 N_A_18 0.00134206f
cc_52 N_NET019_9 N_A_12 0.00842868f
cc_53 N_NET019_8 N_MM11_g 0.0341529f
cc_54 N_NET019_1 N_MM10_g 0.00154355f
cc_55 N_NET019_7 N_B_1 0.00212356f
cc_56 N_NET019_7 N_MM10_g 0.0339634f
cc_57 N_NET019_8 N_NET036_4 0.000422137f
cc_58 N_NET019_7 N_NET036_4 0.000578943f
cc_59 N_NET019_8 N_NET036_1 0.000663427f
cc_60 N_NET019_2 N_MM9_g 0.000904631f
cc_61 N_NET019_8 N_MM9_g 0.034092f
x_PM_XOR2xp5_ASAP7_75t_R%B VSS B N_MM1_g N_MM10_g N_B_1 N_B_6 N_B_7 N_B_5
+ PM_XOR2xp5_ASAP7_75t_R%B
cc_62 N_B_1 N_MM0_g 0.000368993f
cc_63 N_B_6 N_MM0_g 0.000272835f
cc_64 N_B_7 N_MM0_g 0.000327878f
cc_65 N_B_1 N_A_1 0.00179117f
cc_66 N_B_1 N_A_12 0.000424587f
cc_67 N_B_7 N_A_9 0.000482972f
cc_68 N_B_1 N_A_2 0.000487389f
cc_69 N_B_1 N_A_16 0.00196061f
cc_70 N_B_5 N_A_9 0.00216126f
cc_71 N_B_6 N_A_10 0.00485282f
cc_72 N_MM10_g N_MM11_g 0.00490939f
cc_73 N_MM1_g N_MM0_g 0.00743415f
x_PM_XOR2xp5_ASAP7_75t_R%A VSS A N_MM0_g N_MM11_g N_A_1 N_A_12 N_A_9 N_A_2
+ N_A_16 N_A_10 N_A_7 N_A_13 N_A_17 N_A_18 PM_XOR2xp5_ASAP7_75t_R%A
x_PM_XOR2xp5_ASAP7_75t_R%NET036 VSS N_MM9_g N_MM2_s N_MM0_s N_MM1_s N_NET036_14
+ N_NET036_10 N_NET036_4 N_NET036_3 N_NET036_12 N_NET036_1 N_NET036_15
+ N_NET036_16 N_NET036_11 N_NET036_13 N_NET036_18 N_NET036_19
+ PM_XOR2xp5_ASAP7_75t_R%NET036
cc_74 N_NET036_14 N_MM0_g 0.000292027f
cc_75 N_NET036_10 N_A_1 0.000369571f
cc_76 N_NET036_4 N_A_16 0.000498853f
cc_77 N_NET036_3 N_MM0_g 0.000610858f
cc_78 N_NET036_12 N_A_7 0.000769181f
cc_79 N_NET036_4 N_A_12 0.00079663f
cc_80 N_NET036_1 N_A_2 0.00198511f
cc_81 N_NET036_15 N_A_13 0.00162059f
cc_82 N_NET036_4 N_A_10 0.00163508f
cc_83 N_NET036_14 N_A_10 0.00167388f
cc_84 N_NET036_14 N_A_16 0.00260546f
cc_85 N_NET036_16 N_A_13 0.00293113f
cc_86 N_MM9_g N_MM11_g 0.00338312f
cc_87 N_NET036_10 N_MM0_g 0.0263953f
cc_88 N_NET036_11 N_B_7 0.000252713f
cc_89 N_NET036_13 N_B_7 0.000402489f
cc_90 N_NET036_14 N_B_1 0.000724088f
cc_91 N_NET036_4 N_B_5 0.00075426f
cc_92 N_NET036_14 N_B_6 0.000839989f
cc_93 N_NET036_3 N_MM1_g 0.000845936f
cc_94 N_NET036_15 N_B_1 0.000927972f
cc_95 N_NET036_18 N_B_7 0.00264247f
cc_96 N_NET036_4 N_MM1_g 0.00315994f
cc_97 N_NET036_12 N_B_7 0.00328825f
cc_98 N_NET036_10 N_MM1_g 0.0109967f
cc_99 N_NET036_4 N_B_1 0.00488079f
cc_100 N_NET036_14 N_B_5 0.00988383f
cc_101 N_NET036_11 N_MM1_g 0.0500158f
*END of XOR2xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	XNOR2x1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XNOR2x1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XNOR2x1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00618302f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0420733f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0048035f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00655665f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00602407f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00630812f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%NET041 VSS 2 3 1
c1 1 VSS 0.00103441f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5400 $Y2=0.2025
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%NET041__2 VSS 2 3 1
c1 1 VSS 0.00102628f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3240 $Y2=0.2025
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.042214f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%NET43 VSS 2 3 1
c1 1 VSS 0.000993129f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0422992f
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%NET015 VSS 19 41 42 45 46 48 14 2 17 15 1 3 13
+ 16 4
c1 1 VSS 0.00699451f
c2 2 VSS 0.0070312f
c3 3 VSS 0.00711971f
c4 4 VSS 0.00805136f
c5 13 VSS 0.00371853f
c6 14 VSS 0.0033377f
c7 15 VSS 0.00333047f
c8 16 VSS 0.00343456f
c9 17 VSS 0.0334955f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.0675 $X2=0.5920 $Y2=0.0675
r2 48 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.0675 $X2=0.5795 $Y2=0.0675
r3 46 44 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r4 3 44 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r5 15 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r6 45 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r7 42 40 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r8 2 40 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r9 14 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r10 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r11 4 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.0675
+ $X2=0.5940 $Y2=0.0360
r12 3 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r13 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r14 36 37 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.0360 $X2=0.5940 $Y2=0.0360
r15 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5805 $Y2=0.0360
r16 34 35 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.5420
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r17 33 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5240
+ $Y=0.0360 $X2=0.5420 $Y2=0.0360
r18 32 33 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0360 $X2=0.5240 $Y2=0.0360
r19 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4995
+ $Y=0.0360 $X2=0.5130 $Y2=0.0360
r20 30 31 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.4995 $Y2=0.0360
r21 29 30 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r22 28 29 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4430
+ $Y=0.0360 $X2=0.4725 $Y2=0.0360
r23 27 28 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.0360 $X2=0.4430 $Y2=0.0360
r24 26 27 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.4160 $Y2=0.0360
r25 25 26 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r26 24 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3780
+ $Y=0.0360 $X2=0.3915 $Y2=0.0360
r27 23 24 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3670
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r28 22 23 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3440
+ $Y=0.0360 $X2=0.3670 $Y2=0.0360
r29 21 22 10.0272 $w=1.3e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3010
+ $Y=0.0360 $X2=0.3440 $Y2=0.0360
r30 20 21 7.22888 $w=1.3e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3010 $Y2=0.0360
r31 17 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r32 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r33 19 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r34 13 18 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r35 1 13 1e-05
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%Y VSS 31 24 25 50 51 53 55 18 19 4 15 13 1 20 14
+ 16 17 3 2
c1 1 VSS 0.00592342f
c2 2 VSS 0.00286466f
c3 3 VSS 0.00954314f
c4 4 VSS 0.00620283f
c5 13 VSS 0.00202902f
c6 14 VSS 0.00308269f
c7 15 VSS 0.00441579f
c8 16 VSS 0.00260814f
c9 17 VSS 0.0172942f
c10 18 VSS 0.00168787f
c11 19 VSS 0.0137249f
c12 20 VSS 0.000270327f
c13 21 VSS 0.00206731f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5795 $Y=0.2025 $X2=0.5920 $Y2=0.2025
r2 55 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5770 $Y=0.2025 $X2=0.5795 $Y2=0.2025
r3 53 52 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r4 14 52 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r5 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r6 3 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.2025 $X2=0.4465 $Y2=0.2025
r7 15 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r8 50 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r9 4 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5940 $Y=0.2025
+ $X2=0.5940 $Y2=0.2340
r10 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r11 3 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r12 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5805
+ $Y=0.2340 $X2=0.5940 $Y2=0.2340
r13 43 44 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.5510
+ $Y=0.2340 $X2=0.5805 $Y2=0.2340
r14 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.5240
+ $Y=0.2340 $X2=0.5510 $Y2=0.2340
r15 41 42 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.2340 $X2=0.5240 $Y2=0.2340
r16 19 21 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r17 19 41 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.5130 $Y2=0.2340
r18 39 40 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r19 37 40 16.2067 $w=1.3e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4160
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r20 35 36 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r21 17 35 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r22 17 37 1.04935 $w=1.3e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.2340 $X2=0.4160 $Y2=0.2340
r23 21 34 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r24 21 36 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r25 33 34 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1980 $X2=0.4590 $Y2=0.2160
r26 32 33 3.32295 $w=1.3e-08 $l=1.43e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1837 $X2=0.4590 $Y2=0.1980
r27 31 32 1.34084 $w=1.3e-08 $l=5.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4590 $Y2=0.1837
r28 31 30 3.08976 $w=1.3e-08 $l=1.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4590 $Y2=0.1647
r29 29 30 6.58761 $w=1.3e-08 $l=2.82e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1365 $X2=0.4590 $Y2=0.1647
r30 18 28 3.94987 $w=1.50455e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.1080 $X2=0.4590 $Y2=0.0860
r31 18 29 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1080 $X2=0.4590 $Y2=0.1365
r32 27 28 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4455 $Y=0.0860 $X2=0.4590 $Y2=0.0860
r33 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0860 $X2=0.4455 $Y2=0.0860
r34 20 26 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4205
+ $Y=0.0860 $X2=0.4320 $Y2=0.0860
r35 2 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0860
r36 25 23 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r37 2 23 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4320 $Y=0.0675 $X2=0.4465 $Y2=0.0675
r38 13 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r39 24 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r40 1 14 1e-05
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%NET29 VSS 9 10 44 51 52 12 14 1 4 17 13 3 16 11
+ 18 20
c1 1 VSS 0.00580518f
c2 3 VSS 0.0123101f
c3 4 VSS 0.00793166f
c4 9 VSS 0.0434521f
c5 10 VSS 0.0435299f
c6 11 VSS 0.00539043f
c7 12 VSS 0.00778459f
c8 13 VSS 0.0096033f
c9 14 VSS 0.00236428f
c10 15 VSS 0.0016756f
c11 16 VSS 0.00480355f
c12 17 VSS 0.00162915f
c13 18 VSS 0.00145316f
c14 19 VSS 0.0035868f
c15 20 VSS 0.00130373f
r1 52 50 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 3 50 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 51 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1120 $Y2=0.2340
r6 45 46 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r7 13 19 3.94193 $w=1.70327e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1590 $Y=0.2340 $X2=0.1835 $Y2=0.2340
r8 13 46 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r9 11 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r10 44 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r11 4 40 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1750 $Y=0.0675
+ $X2=0.1830 $Y2=0.0960
r12 15 18 2.64331 $w=1.65e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.2160 $X2=0.1835 $Y2=0.1980
r13 15 19 2.23928 $w=1.65e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.2160 $X2=0.1835 $Y2=0.2340
r14 40 41 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.0960 $X2=0.1830 $Y2=0.1130
r15 38 41 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1325 $X2=0.1830 $Y2=0.1130
r16 14 18 6.19173 $w=1.44844e-08 $l=3.1504e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1830 $Y=0.1665 $X2=0.1835 $Y2=0.1980
r17 14 38 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.1665 $X2=0.1830 $Y2=0.1325
r18 18 37 3.27685 $w=1.54359e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1835 $Y=0.1980 $X2=0.2030 $Y2=0.1980
r19 36 37 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2345
+ $Y=0.1980 $X2=0.2030 $Y2=0.1980
r20 35 36 10.7267 $w=1.3e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2805
+ $Y=0.1980 $X2=0.2345 $Y2=0.1980
r21 34 35 12.7088 $w=1.3e-08 $l=5.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3350
+ $Y=0.1980 $X2=0.2805 $Y2=0.1980
r22 16 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3805 $Y=0.1980 $X2=0.4050 $Y2=0.1980
r23 16 34 10.6101 $w=1.3e-08 $l=4.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3805
+ $Y=0.1980 $X2=0.3350 $Y2=0.1980
r24 20 32 5.69636 $w=1.58e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1665
r25 10 29 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r26 17 22 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r27 17 32 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1665
r28 27 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r29 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r30 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r31 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.4145 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r32 22 23 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4145 $Y2=0.1350
r33 1 22 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r34 1 24 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3955
+ $Y=0.1350 $X2=0.3945 $Y2=0.1350
r35 9 22 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r36 9 24 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4050 $Y=0.1350 $X2=0.3945 $Y2=0.1350
r37 9 25 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%A VSS 37 5 6 7 9 1 8 10 11 2 12
c1 1 VSS 0.00705399f
c2 2 VSS 0.00262137f
c3 5 VSS 0.0436343f
c4 6 VSS 0.0435062f
c5 7 VSS 0.0431214f
c6 8 VSS 0.00291781f
c7 9 VSS 0.00478628f
c8 10 VSS 0.00100169f
c9 11 VSS 0.00132692f
c10 12 VSS 0.0389151f
r1 2 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r2 7 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 11 43 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.1980 $X2=0.5670 $Y2=0.1845
r4 11 41 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1980 $X2=0.5670
+ $Y2=0.1890
r5 45 46 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1480
r6 9 43 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1660 $X2=0.5670 $Y2=0.1845
r7 9 46 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1660 $X2=0.5670 $Y2=0.1480
r8 41 43 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.5670 $Y=0.1890 $X2=0.5670
+ $Y2=0.1845
r9 40 41 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M2 $thickness=3.6e-08 $X=0.5425
+ $Y=0.1890 $X2=0.5670 $Y2=0.1890
r10 39 40 30.3147 $w=1.3e-08 $l=1.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.4125
+ $Y=0.1890 $X2=0.5425 $Y2=0.1890
r11 38 39 36.3193 $w=1.3e-08 $l=1.558e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2567 $Y=0.1890 $X2=0.4125 $Y2=0.1890
r12 37 38 9.73567 $w=1.3e-08 $l=4.17e-08 $layer=M2 $thickness=3.6e-08 $X=0.2150
+ $Y=0.1890 $X2=0.2567 $Y2=0.1890
r13 37 36 8.33653 $w=1.3e-08 $l=3.58e-08 $layer=M2 $thickness=3.6e-08 $X=0.2150
+ $Y=0.1890 $X2=0.1792 $Y2=0.1890
r14 35 36 10.3186 $w=1.3e-08 $l=4.42e-08 $layer=M2 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1890 $X2=0.1792 $Y2=0.1890
r15 12 35 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.1235
+ $Y=0.1890 $X2=0.1350 $Y2=0.1890
r16 10 33 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1845
r17 10 35 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1980 $X2=0.1350
+ $Y2=0.1890
r18 33 35 39.0693 $w=9e-09 $l=1.8e-08 $layer=V1 $X=0.1350 $Y=0.1845 $X2=0.1350
+ $Y2=0.1890
r19 32 33 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1620 $X2=0.1350 $Y2=0.1845
r20 30 32 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1435 $X2=0.1350 $Y2=0.1620
r21 29 30 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1435
r22 8 29 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1350
r23 5 24 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r24 24 25 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r25 24 29 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r26 21 25 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1445 $Y2=0.1350
r27 20 21 38.4626 $w=9.3e-09 $l=1.65e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1640 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r28 19 20 58.2767 $w=9.3e-09 $l=2.5e-08 $layer=LIG $thickness=4.8e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1640 $Y2=0.1350
r29 18 19 93.2428 $w=9.3e-09 $l=4e-08 $layer=LIG $thickness=4.8e-08 $X=0.2290
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r30 17 18 95.5738 $w=9.3e-09 $l=4.1e-08 $layer=LIG $thickness=4.8e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2290 $Y2=0.1350
r31 16 17 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r32 6 1 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r33 1 27 7.05813 $w=1.53909e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3080 $Y2=0.1350
r34 6 16 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2970 $Y=0.1350 $X2=0.2845 $Y2=0.1350
r35 6 27 2.64573 $w=2.07209e-07 $l=1.1e-08 $layer=LIG $thickness=5.52727e-08
+ $X=0.2970 $Y=0.1350 $X2=0.3080 $Y2=0.1350
.ends

.subckt PM_XNOR2x1_ASAP7_75t_R%B VSS 34 7 8 9 18 2 10 1 16 13 17 24 11 15 12 3
+ 25 22 14 21 23
c1 1 VSS 0.00882259f
c2 2 VSS 0.00391952f
c3 3 VSS 0.00426351f
c4 7 VSS 0.0818714f
c5 8 VSS 0.0815403f
c6 9 VSS 0.0814524f
c7 10 VSS 0.00855015f
c8 11 VSS 0.0120638f
c9 12 VSS 0.020519f
c10 13 VSS 0.00214248f
c11 14 VSS 0.000361769f
c12 15 VSS 0.000904713f
c13 16 VSS 0.00105789f
c14 17 VSS 0.000401647f
c15 18 VSS 0.00234225f
c16 19 VSS 0.00489083f
c17 20 VSS 0.00201089f
c18 21 VSS 0.00285172f
c19 22 VSS 0.00025296f
c20 23 VSS 0.000639974f
c21 24 VSS 0.000234509f
c22 25 VSS 0.0140309f
r1 2 67 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r2 8 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 3 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
r4 9 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r5 17 67 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3325
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 17 24 2.6649 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3325 $Y=0.1350 $X2=0.3140 $Y2=0.1350
r7 64 65 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1235 $X2=0.5130 $Y2=0.1350
r8 63 64 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1080 $X2=0.5130 $Y2=0.1235
r9 62 63 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0925 $X2=0.5130 $Y2=0.1080
r10 61 62 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0835 $X2=0.5130 $Y2=0.0925
r11 60 61 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0745 $X2=0.5130 $Y2=0.0835
r12 18 60 0.816164 $w=1.3e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.0710 $X2=0.5130 $Y2=0.0745
r13 24 55 1.03257 $w=2.06696e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3140 $Y=0.1350 $X2=0.3140 $Y2=0.1235
r14 58 61 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.5130 $Y=0.0810
+ $X2=0.5130 $Y2=0.0835
r15 57 58 23.2024 $w=1.3e-08 $l=9.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.4135
+ $Y=0.0810 $X2=0.5130 $Y2=0.0810
r16 56 57 23.2024 $w=1.3e-08 $l=9.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0810 $X2=0.4135 $Y2=0.0810
r17 25 56 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M2 $thickness=3.6e-08 $X=0.3015
+ $Y=0.0810 $X2=0.3140 $Y2=0.0810
r18 54 55 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.1080 $X2=0.3140 $Y2=0.1235
r19 53 54 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0925 $X2=0.3140 $Y2=0.1080
r20 16 53 1.16595 $w=1.3e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0875 $X2=0.3140 $Y2=0.0925
r21 16 52 0.991152 $w=1.60769e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.3140 $Y=0.0875 $X2=0.3140 $Y2=0.0810
r22 16 56 70.3248 $w=5e-09 $l=1.8e-08 $layer=V1 $X=0.3140 $Y=0.0875 $X2=0.3140
+ $Y2=0.0810
r23 52 56 27.048 $w=1.3e-08 $l=1.8e-08 $layer=V1 $X=0.3140 $Y=0.0810 $X2=0.3140
+ $Y2=0.0810
r24 50 52 0.663289 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0745 $X2=0.3140 $Y2=0.0810
r25 23 50 0.357156 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0710 $X2=0.3140 $Y2=0.0745
r26 23 51 0.255111 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3140
+ $Y=0.0710 $X2=0.3140 $Y2=0.0685
r27 49 50 5.96826 $w=1.3463e-08 $l=3.35336e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2805 $Y=0.0760 $X2=0.3140 $Y2=0.0745
r28 49 51 5.86622 $w=1.32885e-08 $l=3.43293e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2805 $Y=0.0760 $X2=0.3140 $Y2=0.0685
r29 49 52 6.12133 $w=1.37018e-08 $l=3.38711e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2805 $Y=0.0760 $X2=0.3140 $Y2=0.0810
r30 15 22 3.68021 $w=1.4875e-08 $l=2.15523e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2435 $Y=0.0760 $X2=0.2220 $Y2=0.0745
r31 15 49 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2435
+ $Y=0.0760 $X2=0.2805 $Y2=0.0760
r32 14 21 3.01468 $w=1.741e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2220
+ $Y=0.0560 $X2=0.2220 $Y2=0.0360
r33 14 22 3.33042 $w=1.5027e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2220 $Y=0.0560 $X2=0.2220 $Y2=0.0745
r34 21 47 2.89809 $w=1.53077e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2220 $Y=0.0360 $X2=0.2025 $Y2=0.0360
r35 46 47 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1830
+ $Y=0.0360 $X2=0.2025 $Y2=0.0360
r36 45 46 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.0360 $X2=0.1830 $Y2=0.0360
r37 44 45 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1590 $Y2=0.0360
r38 43 44 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1165
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r39 42 43 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0995
+ $Y=0.0360 $X2=0.1165 $Y2=0.0360
r40 41 42 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0850
+ $Y=0.0360 $X2=0.0995 $Y2=0.0360
r41 12 19 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.0360 $X2=0.0270 $Y2=0.0360
r42 12 41 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.0360 $X2=0.0850 $Y2=0.0360
r43 19 37 4.76361 $w=1.62073e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0635
r44 11 20 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r45 36 37 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1015 $X2=0.0270 $Y2=0.0635
r46 10 20 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1235 $X2=0.0270 $Y2=0.1350
r47 10 36 5.13018 $w=1.3e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1235 $X2=0.0270 $Y2=0.1015
r48 34 13 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r49 13 20 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r50 34 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r51 30 32 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r52 1 29 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r53 1 30 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r54 7 29 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r55 7 30 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends


*
.SUBCKT XNOR2x1_ASAP7_75t_R VSS VDD B A Y
*
* VSS VSS
* VDD VDD
* B B
* A A
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM10@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM11@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM9_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6@2 N_MM6@2_d N_MM9@2_g N_MM6@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5@2 N_MM5@2_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4@2 N_MM4@2_d N_MM10_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM10@2_g N_MM10@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9@2 N_MM9@2_d N_MM9@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XNOR2x1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XNOR2x1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XNOR2x1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_18
cc_1 N_noxref_18_1 N_MM10_g 0.00170667f
cc_2 N_noxref_18_1 N_NET015_16 0.000561092f
cc_3 N_noxref_18_1 N_Y_16 0.0362288f
cc_4 N_noxref_18_1 N_noxref_17_1 0.00179021f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_14
cc_5 N_noxref_14_1 N_A_1 0.00111923f
cc_6 N_noxref_14_1 N_MM2_g 0.00232431f
cc_7 N_noxref_14_1 N_noxref_13_1 0.000901563f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_13
cc_8 N_noxref_13_1 N_A_1 0.000991748f
cc_9 N_noxref_13_1 N_MM2_g 0.00220512f
cc_10 N_noxref_13_1 N_NET29_4 0.00163217f
cc_11 N_noxref_13_1 N_NET29_11 0.0367596f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_16
cc_12 N_noxref_16_1 N_A_1 0.00112832f
cc_13 N_noxref_16_1 N_MM10@2_g 0.00234367f
cc_14 N_noxref_16_1 N_Y_14 0.0354892f
cc_15 N_noxref_16_1 N_noxref_14_1 0.00745617f
cc_16 N_noxref_16_1 N_noxref_15_1 0.000895648f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_15
cc_17 N_noxref_15_1 N_A_1 0.00107765f
cc_18 N_noxref_15_1 N_MM10@2_g 0.00230453f
cc_19 N_noxref_15_1 N_NET29_4 0.00105389f
cc_20 N_noxref_15_1 N_NET015_13 0.0352815f
cc_21 N_noxref_15_1 N_noxref_13_1 0.00729301f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_17
cc_22 N_noxref_17_1 N_MM10_g 0.00163767f
cc_23 N_noxref_17_1 N_NET015_16 0.036104f
cc_24 N_noxref_17_1 N_Y_16 0.000551753f
x_PM_XNOR2x1_ASAP7_75t_R%NET041 VSS N_MM11_d N_MM10_s N_NET041_1
+ PM_XNOR2x1_ASAP7_75t_R%NET041
cc_25 N_NET041_1 N_MM11_g 0.0174109f
cc_26 N_NET041_1 N_MM10_g 0.0173553f
x_PM_XNOR2x1_ASAP7_75t_R%NET041__2 VSS N_MM10@2_s N_MM11@2_d N_NET041__2_1
+ PM_XNOR2x1_ASAP7_75t_R%NET041__2
cc_27 N_NET041__2_1 N_MM11@2_g 0.0172275f
cc_28 N_NET041__2_1 N_MM10@2_g 0.0173927f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_11
cc_29 N_noxref_11_1 N_B_1 0.000239215f
cc_30 N_noxref_11_1 N_MM3_g 0.00229937f
x_PM_XNOR2x1_ASAP7_75t_R%NET43 VSS N_MM3_d N_MM2_s N_NET43_1
+ PM_XNOR2x1_ASAP7_75t_R%NET43
cc_31 N_NET43_1 N_MM3_g 0.0173137f
cc_32 N_NET43_1 N_MM2_g 0.0172255f
x_PM_XNOR2x1_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XNOR2x1_ASAP7_75t_R%noxref_12
cc_33 N_noxref_12_1 N_B_1 0.000238356f
cc_34 N_noxref_12_1 N_MM3_g 0.00222976f
cc_35 N_noxref_12_1 N_noxref_11_1 0.00174589f
x_PM_XNOR2x1_ASAP7_75t_R%NET015 VSS N_MM4_d N_MM5_d N_MM6_s N_MM6@2_s N_MM5@2_d
+ N_MM4@2_d N_NET015_14 N_NET015_2 N_NET015_17 N_NET015_15 N_NET015_1
+ N_NET015_3 N_NET015_13 N_NET015_16 N_NET015_4 PM_XNOR2x1_ASAP7_75t_R%NET015
cc_36 N_NET015_14 N_B_22 0.000130546f
cc_37 N_NET015_14 N_B_18 0.000150005f
cc_38 N_NET015_14 N_B_17 0.000200415f
cc_39 N_NET015_14 N_B_3 0.000231475f
cc_40 N_NET015_14 N_B_16 0.00025862f
cc_41 N_NET015_14 N_B_14 0.000266319f
cc_42 N_NET015_2 N_B_2 0.000288811f
cc_43 N_NET015_17 N_B_16 0.000362069f
cc_44 N_NET015_17 N_B_18 0.000395705f
cc_45 N_NET015_15 N_MM11_g 0.0333679f
cc_46 N_NET015_17 N_B_21 0.00052829f
cc_47 N_NET015_1 N_B_15 0.00164071f
cc_48 N_NET015_14 N_B_2 0.000795625f
cc_49 N_NET015_15 N_B_3 0.00080398f
cc_50 N_NET015_2 N_MM11@2_g 0.00105754f
cc_51 N_NET015_17 N_B_23 0.00106859f
cc_52 N_NET015_3 N_MM11_g 0.00117027f
cc_53 N_NET015_3 N_B_18 0.00180419f
cc_54 N_NET015_17 N_B_15 0.00229649f
cc_55 N_NET015_17 N_B_25 0.00798533f
cc_56 N_NET015_14 N_MM11@2_g 0.0339408f
cc_57 N_NET015_13 N_MM10_g 6.76143e-20
cc_58 N_NET015_13 N_A_12 0.000240667f
cc_59 N_NET015_13 N_A_2 0.000367912f
cc_60 N_NET015_13 N_A_9 0.000457535f
cc_61 N_NET015_16 N_MM10_g 0.0335365f
cc_62 N_NET015_17 N_A_9 0.000504728f
cc_63 N_NET015_16 N_A_2 0.000770932f
cc_64 N_NET015_4 N_MM10_g 0.00118059f
cc_65 N_NET015_1 N_MM10@2_g 0.00150106f
cc_66 N_NET015_13 N_A_1 0.00209001f
cc_67 N_NET015_13 N_MM10@2_g 0.0341815f
cc_68 N_NET015_15 N_MM9_g 0.00043552f
cc_69 N_NET015_13 N_NET29_4 0.000595063f
cc_70 N_NET015_3 N_MM9@2_g 0.000679781f
cc_71 N_NET015_2 N_MM9_g 0.000945238f
cc_72 N_NET015_14 N_NET29_1 0.00141709f
cc_73 N_NET015_14 N_MM9_g 0.0330434f
cc_74 N_NET015_15 N_MM9@2_g 0.0348869f
x_PM_XNOR2x1_ASAP7_75t_R%Y VSS Y N_MM6_d N_MM6@2_d N_MM9_d N_MM9@2_d N_MM10@2_d
+ N_MM10_d N_Y_18 N_Y_19 N_Y_4 N_Y_15 N_Y_13 N_Y_1 N_Y_20 N_Y_14 N_Y_16 N_Y_17
+ N_Y_3 N_Y_2 PM_XNOR2x1_ASAP7_75t_R%Y
cc_75 N_Y_18 N_B_24 8.80943e-20
cc_76 N_Y_18 N_MM11_g 8.83417e-20
cc_77 N_Y_18 N_B_2 0.000207543f
cc_78 N_Y_18 N_MM11@2_g 9.56377e-20
cc_79 N_Y_18 N_B_17 0.000315935f
cc_80 N_Y_19 N_B_18 0.000189844f
cc_81 N_Y_4 N_MM11_g 0.000195503f
cc_82 N_Y_15 N_B_3 0.00021819f
cc_83 N_Y_13 N_MM11_g 0.000310666f
cc_84 N_Y_1 N_MM11@2_g 0.000327164f
cc_85 N_Y_13 N_MM11@2_g 0.000332724f
cc_86 N_Y_18 N_B_3 0.000360359f
cc_87 N_Y_20 N_B_18 0.00062259f
cc_88 N_Y_20 N_B_25 0.00194486f
cc_89 N_Y_18 N_B_18 0.00408482f
cc_90 N_Y_14 N_A_12 0.000119571f
cc_91 N_Y_14 N_A_9 0.000258271f
cc_92 N_Y_14 N_A_11 0.000293883f
cc_93 N_Y_14 N_A_2 0.000341722f
cc_94 N_Y_16 N_MM10_g 0.0342858f
cc_95 N_Y_4 N_A_9 0.000789195f
cc_96 N_Y_16 N_A_2 0.000841848f
cc_97 N_Y_18 N_A_12 0.00127518f
cc_98 N_Y_1 N_MM10@2_g 0.00178994f
cc_99 N_Y_4 N_MM10_g 0.00196255f
cc_100 N_Y_14 N_A_1 0.00234655f
cc_101 N_Y_17 N_A_12 0.00430251f
cc_102 N_Y_19 N_A_11 0.00674368f
cc_103 N_Y_14 N_MM10@2_g 0.0348722f
cc_104 N_Y_20 N_NET29_17 0.000547973f
cc_105 N_Y_3 N_NET29_1 0.000600151f
cc_106 N_Y_15 N_MM9_g 0.0305377f
cc_107 N_Y_1 N_NET29_16 0.00112339f
cc_108 N_Y_17 N_NET29_20 0.00152135f
cc_109 N_Y_2 N_MM9_g 0.00171566f
cc_110 N_Y_3 N_MM9_g 0.00212767f
cc_111 N_Y_18 N_NET29_17 0.00414763f
cc_112 N_Y_15 N_NET29_1 0.00506041f
cc_113 N_Y_17 N_NET29_16 0.0119616f
cc_114 N_Y_13 N_MM9@2_g 0.0367148f
cc_115 N_Y_13 N_MM9_g 0.0684685f
cc_116 N_Y_18 N_NET015_3 0.000288153f
cc_117 N_Y_13 N_NET015_14 0.00168914f
cc_118 N_Y_13 N_NET015_15 0.000562833f
cc_119 N_Y_2 N_NET015_17 0.000686504f
cc_120 N_Y_2 N_NET015_3 0.00163244f
cc_121 N_Y_20 N_NET015_17 0.00366143f
cc_122 N_Y_2 N_NET015_2 0.00594775f
x_PM_XNOR2x1_ASAP7_75t_R%NET29 VSS N_MM9_g N_MM9@2_g N_MM2_d N_MM1_d N_MM0_d
+ N_NET29_12 N_NET29_14 N_NET29_1 N_NET29_4 N_NET29_17 N_NET29_13 N_NET29_3
+ N_NET29_16 N_NET29_11 N_NET29_18 N_NET29_20 PM_XNOR2x1_ASAP7_75t_R%NET29
cc_123 N_NET29_12 N_B_3 0.000134467f
cc_124 N_NET29_12 N_B_1 0.00107704f
cc_125 N_NET29_12 N_B_13 0.000200342f
cc_126 N_NET29_12 N_B_16 0.000216423f
cc_127 N_NET29_14 N_B_14 0.000350978f
cc_128 N_NET29_1 N_B_17 0.000361095f
cc_129 N_NET29_4 N_B_22 0.000374307f
cc_130 N_NET29_1 N_B_3 0.000375819f
cc_131 N_NET29_14 N_B_15 0.000517096f
cc_132 N_NET29_17 N_B_25 0.000553477f
cc_133 N_NET29_1 N_B_2 0.00209108f
cc_134 N_NET29_13 N_B_11 0.000711692f
cc_135 N_NET29_3 N_MM3_g 0.000976626f
cc_136 N_NET29_16 N_B_24 0.00216164f
cc_137 N_NET29_17 N_B_17 0.00253321f
cc_138 N_NET29_14 N_B_22 0.00301709f
cc_139 N_MM9@2_g N_MM11_g 0.00336438f
cc_140 N_MM9_g N_MM11@2_g 0.00341604f
cc_141 N_NET29_4 N_B_12 0.00386859f
cc_142 N_NET29_12 N_MM3_g 0.0356241f
cc_143 N_NET29_11 N_MM10@2_g 0.000151625f
cc_144 N_NET29_11 N_A_10 0.000784371f
cc_145 N_NET29_11 N_A_12 0.000281972f
cc_146 N_NET29_12 N_MM2_g 0.0156917f
cc_147 N_NET29_13 N_A_8 0.000449921f
cc_148 N_NET29_4 N_A_1 0.00572061f
cc_149 N_NET29_17 N_A_12 0.00065612f
cc_150 N_NET29_18 N_A_10 0.000750737f
cc_151 N_NET29_3 N_A_1 0.000834757f
cc_152 N_NET29_3 N_MM2_g 0.00144526f
cc_153 N_NET29_4 N_MM2_g 0.00289879f
cc_154 N_NET29_13 N_A_10 0.00493164f
cc_155 N_NET29_14 N_A_8 0.00580697f
cc_156 N_NET29_16 N_A_12 0.00758542f
cc_157 N_NET29_11 N_MM2_g 0.0548322f
x_PM_XNOR2x1_ASAP7_75t_R%A VSS A N_MM2_g N_MM10@2_g N_MM10_g N_A_9 N_A_1 N_A_8
+ N_A_10 N_A_11 N_A_2 N_A_12 PM_XNOR2x1_ASAP7_75t_R%A
cc_158 N_A_9 N_MM3_g 7.3618e-20
cc_159 N_A_1 N_MM3_g 0.00010486f
cc_160 N_A_8 N_MM3_g 0.000113357f
cc_161 N_A_9 N_B_18 0.00319957f
cc_162 N_A_1 N_B_2 0.000653227f
cc_163 N_A_8 N_B_10 0.000242425f
cc_164 N_A_1 N_B_1 0.0014196f
cc_165 N_A_1 N_B_16 0.000357919f
cc_166 N_A_10 N_B_13 0.000371067f
cc_167 N_A_1 N_B_17 0.000396773f
cc_168 N_A_11 N_B_18 0.000422964f
cc_169 N_A_1 N_B_24 0.00044829f
cc_170 N_A_10 N_B_11 0.000471084f
cc_171 N_A_1 N_B_15 0.000493497f
cc_172 N_A_8 N_B_12 0.000615838f
cc_173 N_A_2 N_B_3 0.00224312f
cc_174 N_A_8 N_B_13 0.00175969f
cc_175 N_A_12 N_B_25 0.00217005f
cc_176 N_A_1 N_B_22 0.00225076f
cc_177 N_A_12 N_B_17 0.00403854f
cc_178 N_MM10@2_g N_MM11@2_g 0.00492342f
cc_179 N_MM10_g N_MM11_g 0.00498308f
cc_180 N_MM2_g N_MM3_g 0.00527778f
x_PM_XNOR2x1_ASAP7_75t_R%B VSS B N_MM3_g N_MM11@2_g N_MM11_g N_B_18 N_B_2
+ N_B_10 N_B_1 N_B_16 N_B_13 N_B_17 N_B_24 N_B_11 N_B_15 N_B_12 N_B_3 N_B_25
+ N_B_22 N_B_14 N_B_21 N_B_23 PM_XNOR2x1_ASAP7_75t_R%B
*END of XNOR2x1_ASAP7_75t_R.pxi
.ENDS
** Design:	XNOR2x2_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XNOR2x2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XNOR2x2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XNOR2x2_ASAP7_75t_R%NET048 VSS 2 3 1
c1 1 VSS 0.000947286f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3780 $Y2=0.2025
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%NET047 VSS 2 3 1
c1 1 VSS 0.00103195f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00470703f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00612269f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00485201f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00495025f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0422921f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.00452996f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%NET019 VSS 12 13 19 7 8 1 9 2
c1 1 VSS 0.00722442f
c2 2 VSS 0.00755597f
c3 7 VSS 0.003403f
c4 8 VSS 0.00371027f
c5 9 VSS 0.0132417f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2140 $Y2=0.2025
r2 19 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r3 2 16 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.2340
r4 15 16 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1665
+ $Y=0.2340 $X2=0.2160 $Y2=0.2340
r5 14 15 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.2340 $X2=0.1665 $Y2=0.2340
r6 9 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r7 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r8 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r9 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r10 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r11 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0310723f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.0422851f
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%Y VSS 21 16 17 28 29 10 7 8 9 11 1 2
c1 1 VSS 0.00996353f
c2 2 VSS 0.0104537f
c3 7 VSS 0.00449025f
c4 8 VSS 0.00447206f
c5 9 VSS 0.00868712f
c6 10 VSS 0.00842493f
c7 11 VSS 0.00702617f
c8 12 VSS 0.00336381f
c9 13 VSS 0.00344625f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 28 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r6 10 13 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5265 $Y=0.2340 $X2=0.5670 $Y2=0.2340
r7 10 24 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.5265
+ $Y=0.2340 $X2=0.4860 $Y2=0.2340
r8 13 23 9.07762 $w=1.49174e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.2340 $X2=0.5670 $Y2=0.1880
r9 22 23 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1495 $X2=0.5670 $Y2=0.1880
r10 21 22 0.46638 $w=1.3e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1475 $X2=0.5670 $Y2=0.1495
r11 21 20 9.91057 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1475 $X2=0.5670 $Y2=0.1050
r12 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0540 $X2=0.5670 $Y2=0.0360
r13 11 20 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0540 $X2=0.5670 $Y2=0.1050
r14 12 19 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5670 $Y=0.0360 $X2=0.5265 $Y2=0.0360
r15 18 19 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0360 $X2=0.5265 $Y2=0.0360
r16 9 18 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4745
+ $Y=0.0360 $X2=0.4860 $Y2=0.0360
r17 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r18 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r19 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r20 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r21 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%B VSS 20 3 4 5 1 6
c1 1 VSS 0.0094723f
c2 3 VSS 0.0466241f
c3 4 VSS 0.0358912f
c4 5 VSS 0.00391138f
c5 6 VSS 0.00393377f
r1 6 23 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1980 $X2=0.3510 $Y2=0.1665
r2 3 17 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r3 21 23 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1435 $X2=0.3510 $Y2=0.1665
r4 20 21 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1435
r5 20 5 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1265
r6 15 17 10.5547 $w=1.466e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r7 14 15 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2015 $Y2=0.1350
r8 13 14 96.7394 $w=9.3e-09 $l=4.15e-08 $layer=LIG $thickness=4.8e-08 $X=0.2575
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r9 12 13 97.9049 $w=9.3e-09 $l=4.2e-08 $layer=LIG $thickness=4.8e-08 $X=0.2995
+ $Y=0.1350 $X2=0.2575 $Y2=0.1350
r10 11 12 57.1112 $w=9.3e-09 $l=2.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.2995 $Y2=0.1350
r11 10 11 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r12 9 19 1.40189 $w=1.265e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.3605
+ $Y=0.1350 $X2=0.3615 $Y2=0.1350
r13 8 9 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3605 $Y2=0.1350
r14 20 8 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r15 1 8 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.3415
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r16 1 10 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3415 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r17 4 8 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r18 4 10 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r19 4 19 1.4802 $w=2.16633e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3615 $Y2=0.1350
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%NET036 VSS 9 39 42 43 3 4 14 15 1 13 12 10 11 17
+ 16
c1 1 VSS 0.0018661f
c2 3 VSS 0.00615017f
c3 4 VSS 0.00760803f
c4 9 VSS 0.0422063f
c5 10 VSS 0.00585306f
c6 11 VSS 0.00466475f
c7 12 VSS 0.00166972f
c8 13 VSS 0.00542662f
c9 14 VSS 0.00183437f
c10 15 VSS 0.00185258f
c11 16 VSS 0.000463261f
c12 17 VSS 0.000492684f
r1 43 41 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0540 $X2=0.3925 $Y2=0.0540
r2 4 41 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0540 $X2=0.3925 $Y2=0.0540
r3 10 4 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0540 $X2=0.3780 $Y2=0.0540
r4 42 10 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0540 $X2=0.3635 $Y2=0.0540
r5 39 38 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r6 11 38 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3260 $Y=0.2025 $X2=0.3385 $Y2=0.2025
r7 4 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0540
+ $X2=0.3745 $Y2=0.0720
r8 3 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3115 $Y=0.2025
+ $X2=0.3110 $Y2=0.1770
r9 32 33 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0720 $X2=0.3745 $Y2=0.0720
r10 31 32 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.0720 $X2=0.3645 $Y2=0.0720
r11 15 17 3.48349 $w=1.525e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.0720 $X2=0.3110 $Y2=0.0720
r12 15 31 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.0720 $X2=0.3510 $Y2=0.0720
r13 27 28 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.1455 $X2=0.3110 $Y2=0.1770
r14 26 27 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.1135 $X2=0.3110 $Y2=0.1455
r15 14 17 3.94987 $w=1.50455e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3110 $Y=0.0940 $X2=0.3110 $Y2=0.0720
r16 14 26 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.0940 $X2=0.3110 $Y2=0.1135
r17 17 25 3.60008 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3110 $Y=0.0720 $X2=0.2905 $Y2=0.0720
r18 24 25 18.422 $w=1.3e-08 $l=7.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2115
+ $Y=0.0720 $X2=0.2905 $Y2=0.0720
r19 23 24 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0720 $X2=0.2115 $Y2=0.0720
r20 22 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1125
+ $Y=0.0720 $X2=0.1350 $Y2=0.0720
r21 13 16 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0945 $Y=0.0720 $X2=0.0810 $Y2=0.0720
r22 13 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0720 $X2=0.1125 $Y2=0.0720
r23 16 21 4.9968 $w=1.60947e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0720 $X2=0.0810 $Y2=0.1005
r24 12 19 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1230 $X2=0.0810 $Y2=0.1350
r25 12 21 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1230 $X2=0.0810 $Y2=0.1005
r26 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r27 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r28 3 11 1e-05
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%A VSS 26 5 6 13 2 9 8 15 1 7 10 11 12 16
c1 1 VSS 0.00548541f
c2 2 VSS 0.00597406f
c3 5 VSS 0.082493f
c4 6 VSS 0.0826653f
c5 7 VSS 0.00198108f
c6 8 VSS 0.00326606f
c7 9 VSS 0.00127069f
c8 10 VSS 0.0141881f
c9 11 VSS 0.00361298f
c10 12 VSS 0.00132042f
c11 13 VSS 0.00107122f
c12 14 VSS 0.00298572f
c13 15 VSS 0.00176414f
c14 16 VSS 0.00343441f
r1 1 39 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r2 5 1 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 39 40 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1465
r4 7 12 4.41382 $w=1.63923e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1660 $X2=0.1350 $Y2=0.1920
r5 7 40 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1660 $X2=0.1350 $Y2=0.1465
r6 12 37 10.4768 $w=1.38654e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1920 $X2=0.1870 $Y2=0.1920
r7 8 13 3.92057 $w=1.38108e-08 $l=2.5224e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2455 $Y=0.1920 $X2=0.2700 $Y2=0.1980
r8 8 37 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2455
+ $Y=0.1920 $X2=0.1870 $Y2=0.1920
r9 13 35 1.0057 $w=1.55e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.1980 $X2=0.2700 $Y2=0.2040
r10 9 14 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2160 $X2=0.2700 $Y2=0.2340
r11 9 35 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2160 $X2=0.2700 $Y2=0.2040
r12 14 34 3.13128 $w=1.51951e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2700 $Y=0.2340 $X2=0.2905 $Y2=0.2340
r13 33 34 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.3110
+ $Y=0.2340 $X2=0.2905 $Y2=0.2340
r14 32 33 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3310
+ $Y=0.2340 $X2=0.3110 $Y2=0.2340
r15 31 32 6.99569 $w=1.3e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.3610
+ $Y=0.2340 $X2=0.3310 $Y2=0.2340
r16 30 31 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3855
+ $Y=0.2340 $X2=0.3610 $Y2=0.2340
r17 10 16 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4065 $Y=0.2340 $X2=0.4310 $Y2=0.2340
r18 10 30 4.89699 $w=1.3e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4065
+ $Y=0.2340 $X2=0.3855 $Y2=0.2340
r19 16 29 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.2340 $X2=0.4310 $Y2=0.2160
r20 28 29 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1980 $X2=0.4310 $Y2=0.2160
r21 27 28 4.4889 $w=1.3e-08 $l=1.93e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1787 $X2=0.4310 $Y2=0.1980
r22 26 27 2.50679 $w=1.3e-08 $l=1.07e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1680 $X2=0.4310 $Y2=0.1787
r23 26 25 2.04041 $w=1.3e-08 $l=8.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1680 $X2=0.4310 $Y2=0.1592
r24 11 23 0.867186 $w=1.3625e-08 $l=1.51162e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4310 $Y=0.1475 $X2=0.4225 $Y2=0.1350
r25 11 25 2.73998 $w=1.3e-08 $l=1.17e-08 $layer=M1 $thickness=3.6e-08 $X=0.4310
+ $Y=0.1475 $X2=0.4310 $Y2=0.1592
r26 22 23 0.983781 $w=1.35556e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.4180 $Y=0.1350 $X2=0.4225 $Y2=0.1350
r27 21 22 3.03147 $w=1.3e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4180 $Y2=0.1350
r28 20 21 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3940
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r29 15 20 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1350 $X2=0.3940 $Y2=0.1350
r30 6 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r31 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends

.subckt PM_XNOR2x2_ASAP7_75t_R%XOR VSS 12 13 49 54 58 15 3 19 18 5 16 25 4 17
+ 14 23 1 20 21 26 24
c1 1 VSS 0.00710959f
c2 3 VSS 0.00813516f
c3 4 VSS 0.00573398f
c4 5 VSS 0.00574939f
c5 12 VSS 0.0803064f
c6 13 VSS 0.0808523f
c7 14 VSS 0.00582718f
c8 15 VSS 0.00502677f
c9 16 VSS 0.00458646f
c10 17 VSS 0.0075343f
c11 18 VSS 0.03657f
c12 19 VSS 0.000698228f
c13 20 VSS 0.00119194f
c14 21 VSS 0.0020421f
c15 22 VSS 0.00341428f
c16 23 VSS 0.00658069f
c17 24 VSS 0.00300792f
c18 25 VSS 0.000815473f
c19 26 VSS 0.000465095f
r1 58 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 16 57 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 4 56 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 55 56 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 23 52 3.71668 $w=1.51429e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2130
r6 23 55 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 54 53 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r8 14 53 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r9 51 52 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1750 $X2=0.0270 $Y2=0.2130
r10 50 51 16.0901 $w=1.3e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1060 $X2=0.0270 $Y2=0.1750
r11 17 22 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.0360
r12 17 50 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0540 $X2=0.0270 $Y2=0.1060
r13 15 5 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2140 $Y2=0.0675
r14 49 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r15 3 45 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r16 22 44 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r17 5 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0540
+ $X2=0.2160 $Y2=0.0360
r18 44 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r19 43 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r20 41 42 21.5701 $w=1.3e-08 $l=9.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.3085 $Y2=0.0360
r21 40 41 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.1395
+ $Y=0.0360 $X2=0.2160 $Y2=0.0360
r22 40 43 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.1395
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r23 18 24 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4075 $Y=0.0360 $X2=0.4320 $Y2=0.0360
r24 18 42 23.0858 $w=1.3e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4075
+ $Y=0.0360 $X2=0.3085 $Y2=0.0360
r25 19 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0540 $X2=0.4320 $Y2=0.0720
r26 19 24 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0540 $X2=0.4320 $Y2=0.0360
r27 25 39 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4320 $Y=0.0720 $X2=0.4565 $Y2=0.0720
r28 20 26 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4745 $Y=0.0720 $X2=0.4860 $Y2=0.0720
r29 20 39 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4745
+ $Y=0.0720 $X2=0.4565 $Y2=0.0720
r30 26 36 3.48106 $w=1.70091e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.0720 $X2=0.4860 $Y2=0.0940
r31 13 33 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r32 35 36 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1165 $X2=0.4860 $Y2=0.0940
r33 21 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4860 $Y=0.1350
+ $X2=0.4860 $Y2=0.1350
r34 21 35 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.1350 $X2=0.4860 $Y2=0.1165
r35 31 33 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.5005 $Y=0.1350 $X2=0.5130 $Y2=0.1350
r36 30 31 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4860 $Y=0.1350 $X2=0.5005 $Y2=0.1350
r37 29 30 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4715 $Y=0.1350 $X2=0.4860 $Y2=0.1350
r38 12 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r39 1 28 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4485 $Y2=0.1350
r40 1 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r41 12 28 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.4590 $Y=0.1350 $X2=0.4485 $Y2=0.1350
r42 12 29 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.4590 $Y=0.1350 $X2=0.4715 $Y2=0.1350
r43 4 16 1e-05
r44 3 14 1e-05
.ends


*
.SUBCKT XNOR2x2_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM9 VSS N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VSS N_MM11_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM10_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 VSS N_MM2_g N_MM1_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM0 VSS N_MM3_g N_MM0_s VSS nmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM13 VSS N_MM12_g N_MM13_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13@2 VSS N_MM12@2_g N_MM13@2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM9_g N_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 VDD N_MM11_g N_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 VDD N_MM10_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 VDD N_MM3_g N_MM3_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 VDD N_MM12_g N_MM12_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12@2 VDD N_MM12@2_g N_MM12@2_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XNOR2x2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XNOR2x2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XNOR2x2_ASAP7_75t_R%NET048 VSS N_MM2_d N_MM3_s N_NET048_1
+ PM_XNOR2x2_ASAP7_75t_R%NET048
cc_1 N_NET048_1 N_MM3_g 0.0173106f
cc_2 N_NET048_1 N_MM2_g 0.0174492f
x_PM_XNOR2x2_ASAP7_75t_R%NET047 VSS N_MM11_s N_MM10_d N_NET047_1
+ PM_XNOR2x2_ASAP7_75t_R%NET047
cc_3 N_NET047_1 N_MM11_g 0.0173114f
cc_4 N_NET047_1 N_MM10_g 0.0173033f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_16
cc_5 N_noxref_16_1 N_NET036_3 0.00158325f
cc_6 N_noxref_16_1 N_NET036_11 0.0366845f
cc_7 N_noxref_16_1 N_B_1 0.00100322f
cc_8 N_noxref_16_1 N_MM2_g 0.00228811f
cc_9 N_noxref_16_1 N_noxref_14_1 0.00730784f
cc_10 N_noxref_16_1 N_noxref_15_1 0.000968181f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_14
cc_11 N_noxref_14_1 N_NET036_3 0.0010071f
cc_12 N_noxref_14_1 N_B_1 0.00108511f
cc_13 N_noxref_14_1 N_MM10_g 0.00229947f
cc_14 N_noxref_14_1 N_NET019_8 0.0352254f
cc_15 N_noxref_14_1 N_noxref_13_1 0.000896035f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_12
cc_16 N_noxref_12_1 N_MM9_g 0.00145195f
cc_17 N_noxref_12_1 N_XOR_17 0.000326924f
cc_18 N_noxref_12_1 N_XOR_4 0.000509729f
cc_19 N_noxref_12_1 N_XOR_16 0.0375221f
cc_20 N_noxref_12_1 N_noxref_11_1 0.00176442f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_13
cc_21 N_noxref_13_1 N_B_1 0.00114472f
cc_22 N_noxref_13_1 N_MM10_g 0.00235887f
cc_23 N_noxref_13_1 N_XOR_15 0.0370192f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_17
cc_24 N_noxref_17_1 N_MM12@2_g 0.00148142f
cc_25 N_noxref_17_1 N_Y_7 0.000828717f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_11
cc_26 N_noxref_11_1 N_MM9_g 0.0014537f
cc_27 N_noxref_11_1 N_XOR_17 0.000325763f
cc_28 N_noxref_11_1 N_XOR_3 0.000508146f
cc_29 N_noxref_11_1 N_XOR_14 0.0377831f
x_PM_XNOR2x2_ASAP7_75t_R%NET019 VSS N_MM6_d N_MM4_s N_MM5_s N_NET019_7
+ N_NET019_8 N_NET019_1 N_NET019_9 N_NET019_2 PM_XNOR2x2_ASAP7_75t_R%NET019
cc_30 N_NET019_7 N_NET036_3 0.000413152f
cc_31 N_NET019_8 N_NET036_3 0.000569255f
cc_32 N_NET019_7 N_NET036_1 0.000633317f
cc_33 N_NET019_1 N_MM9_g 0.000880437f
cc_34 N_NET019_7 N_MM9_g 0.0343657f
cc_35 N_NET019_7 N_A_8 0.000405388f
cc_36 N_NET019_1 N_A_7 0.000505198f
cc_37 N_NET019_7 N_A_1 0.00073898f
cc_38 N_NET019_9 N_A_12 0.000949923f
cc_39 N_NET019_2 N_A_8 0.00106805f
cc_40 N_NET019_1 N_MM11_g 0.00124476f
cc_41 N_NET019_9 N_A_8 0.00718295f
cc_42 N_NET019_7 N_MM11_g 0.0347456f
cc_43 N_NET019_2 N_MM10_g 0.00153066f
cc_44 N_NET019_8 N_B_1 0.00218126f
cc_45 N_NET019_8 N_MM10_g 0.0339542f
cc_46 N_NET019_1 N_XOR_16 0.00112738f
cc_47 N_NET019_9 N_XOR_23 0.000886396f
cc_48 N_NET019_1 N_XOR_4 0.00404768f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_15
cc_49 N_noxref_15_1 N_NET036_10 0.000487659f
cc_50 N_noxref_15_1 N_B_1 0.00141509f
cc_51 N_noxref_15_1 N_MM2_g 0.00431058f
cc_52 N_noxref_15_1 N_XOR_15 0.000553208f
cc_53 N_noxref_15_1 N_noxref_13_1 0.0075103f
x_PM_XNOR2x2_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1
+ PM_XNOR2x2_ASAP7_75t_R%noxref_18
cc_54 N_noxref_18_1 N_MM12@2_g 0.00147039f
cc_55 N_noxref_18_1 N_Y_8 0.000835873f
cc_56 N_noxref_18_1 N_noxref_17_1 0.00176783f
x_PM_XNOR2x2_ASAP7_75t_R%Y VSS Y N_MM13_s N_MM13@2_s N_MM12_s N_MM12@2_s N_Y_10
+ N_Y_7 N_Y_8 N_Y_9 N_Y_11 N_Y_1 N_Y_2 PM_XNOR2x2_ASAP7_75t_R%Y
cc_57 N_Y_10 N_A_11 0.000911626f
cc_58 N_Y_10 N_A_16 0.00238052f
cc_59 N_Y_7 N_XOR_21 0.000297506f
cc_60 N_Y_7 N_XOR_26 0.000368001f
cc_61 N_Y_7 N_XOR_24 0.000384399f
cc_62 N_Y_7 N_XOR_1 0.000736222f
cc_63 N_Y_8 N_MM12_g 0.0307388f
cc_64 N_Y_9 N_XOR_20 0.00096761f
cc_65 N_Y_11 N_XOR_1 0.00129482f
cc_66 N_Y_1 N_XOR_21 0.00173713f
cc_67 N_Y_2 N_MM12_g 0.00197319f
cc_68 N_Y_1 N_MM12_g 0.00265113f
cc_69 N_Y_9 N_XOR_26 0.00327699f
cc_70 N_Y_8 N_XOR_1 0.00424172f
cc_71 N_Y_7 N_MM12@2_g 0.0370791f
cc_72 N_Y_7 N_MM12_g 0.0683314f
x_PM_XNOR2x2_ASAP7_75t_R%B VSS B N_MM10_g N_MM2_g N_B_5 N_B_1 N_B_6
+ PM_XNOR2x2_ASAP7_75t_R%B
cc_73 N_B_5 N_NET036_11 0.000294781f
cc_74 N_MM2_g N_NET036_4 0.000578459f
cc_75 N_B_5 N_NET036_3 0.000641817f
cc_76 N_B_1 N_NET036_13 0.000774613f
cc_77 N_B_6 N_NET036_14 0.000807778f
cc_78 N_B_1 N_NET036_14 0.000857216f
cc_79 N_B_5 N_NET036_15 0.00108637f
cc_80 N_MM2_g N_NET036_3 0.00321465f
cc_81 N_MM2_g N_NET036_10 0.0109107f
cc_82 N_B_1 N_NET036_3 0.00511453f
cc_83 N_B_5 N_NET036_14 0.00809403f
cc_84 N_MM2_g N_NET036_11 0.0498773f
cc_85 N_B_1 N_MM3_g 0.00113007f
cc_86 N_B_1 N_A_1 0.000480419f
cc_87 N_B_1 N_A_2 0.00135654f
cc_88 N_B_6 N_A_11 0.000647259f
cc_89 N_B_1 N_A_13 0.00203722f
cc_90 N_B_5 N_A_15 0.00255979f
cc_91 N_MM10_g N_MM11_g 0.00490625f
cc_92 N_B_6 N_A_10 0.00507159f
cc_93 N_MM2_g N_MM3_g 0.00753318f
x_PM_XNOR2x2_ASAP7_75t_R%NET036 VSS N_MM9_g N_MM2_s N_MM1_s N_MM0_s N_NET036_3
+ N_NET036_4 N_NET036_14 N_NET036_15 N_NET036_1 N_NET036_13 N_NET036_12
+ N_NET036_10 N_NET036_11 N_NET036_17 N_NET036_16 PM_XNOR2x2_ASAP7_75t_R%NET036
x_PM_XNOR2x2_ASAP7_75t_R%A VSS A N_MM11_g N_MM3_g N_A_13 N_A_2 N_A_9 N_A_8
+ N_A_15 N_A_1 N_A_7 N_A_10 N_A_11 N_A_12 N_A_16 PM_XNOR2x2_ASAP7_75t_R%A
cc_94 N_A_13 N_NET036_3 0.000358005f
cc_95 N_A_2 N_NET036_4 0.000387185f
cc_96 N_A_9 N_NET036_14 0.00044886f
cc_97 N_MM3_g N_NET036_4 0.00051223f
cc_98 N_A_8 N_NET036_3 0.000873352f
cc_99 N_A_15 N_NET036_15 0.00090191f
cc_100 N_A_1 N_NET036_1 0.00192212f
cc_101 N_A_7 N_NET036_13 0.00156287f
cc_102 N_A_10 N_NET036_3 0.00162945f
cc_103 N_A_10 N_NET036_14 0.00164091f
cc_104 N_A_7 N_NET036_12 0.00285703f
cc_105 N_A_13 N_NET036_14 0.00307169f
cc_106 N_MM11_g N_MM9_g 0.00336305f
cc_107 N_MM3_g N_NET036_10 0.0260557f
x_PM_XNOR2x2_ASAP7_75t_R%XOR VSS N_MM12_g N_MM12@2_g N_MM10_s N_MM9_s N_MM6_s
+ N_XOR_15 N_XOR_3 N_XOR_19 N_XOR_18 N_XOR_5 N_XOR_16 N_XOR_25 N_XOR_4 N_XOR_17
+ N_XOR_14 N_XOR_23 N_XOR_1 N_XOR_20 N_XOR_21 N_XOR_26 N_XOR_24
+ PM_XNOR2x2_ASAP7_75t_R%XOR
cc_108 N_XOR_15 N_MM9_g 9.16273e-20
cc_109 N_XOR_3 N_MM9_g 0.00158853f
cc_110 N_XOR_19 N_MM9_g 0.000209293f
cc_111 N_XOR_18 N_NET036_14 0.000287674f
cc_112 N_XOR_5 N_NET036_13 0.00154128f
cc_113 N_XOR_16 N_MM9_g 0.0156007f
cc_114 N_XOR_18 N_NET036_4 0.000979762f
cc_115 N_XOR_25 N_NET036_15 0.000487566f
cc_116 N_XOR_3 N_NET036_1 0.000911857f
cc_117 N_XOR_4 N_MM9_g 0.00106956f
cc_118 N_XOR_18 N_NET036_17 0.00117243f
cc_119 N_XOR_16 N_NET036_1 0.00163646f
cc_120 N_XOR_18 N_NET036_16 0.00172118f
cc_121 N_XOR_18 N_NET036_15 0.00299584f
cc_122 N_XOR_17 N_NET036_12 0.00469108f
cc_123 N_XOR_18 N_NET036_13 0.021247f
cc_124 N_XOR_14 N_MM9_g 0.054457f
cc_125 N_XOR_15 N_MM3_g 9.59848e-20
cc_126 N_XOR_3 N_MM3_g 0.000110053f
cc_127 N_XOR_16 N_MM3_g 0.0001143f
cc_128 N_XOR_5 N_MM3_g 0.000209786f
cc_129 N_XOR_23 N_MM3_g 0.000229502f
cc_130 N_XOR_1 N_MM3_g 0.000247797f
cc_131 N_XOR_1 N_A_2 0.00133411f
cc_132 N_XOR_20 N_A_15 0.000264297f
cc_133 N_XOR_17 N_A_7 0.000268729f
cc_134 N_XOR_5 N_MM11_g 0.000305078f
cc_135 N_XOR_18 N_A_7 0.000314587f
cc_136 N_XOR_14 N_MM11_g 0.000342637f
cc_137 N_XOR_4 N_A_7 0.000370581f
cc_138 N_XOR_25 N_A_15 0.000827687f
cc_139 N_XOR_21 N_A_11 0.000834709f
cc_140 N_XOR_21 N_A_15 0.00187171f
cc_141 N_MM12_g N_MM3_g 0.00385091f
cc_142 N_XOR_25 N_B_5 0.000201468f
cc_143 N_XOR_5 N_MM10_g 0.00180505f
cc_144 N_XOR_15 N_B_1 0.00246742f
cc_145 N_XOR_15 N_MM10_g 0.0365167f
*END of XNOR2x2_ASAP7_75t_R.pxi
.ENDS
** Design:	XNOR2xp5_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "XNOR2xp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "XNOR2xp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00550289f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00461933f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0315449f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00619159f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00493991f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.00485709f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%Y VSS 22 18 31 33 1 11 12 3 2 13 10 14 15
c1 1 VSS 0.00656948f
c2 2 VSS 0.00602502f
c3 3 VSS 0.00787229f
c4 10 VSS 0.0026745f
c5 11 VSS 0.00343129f
c6 12 VSS 0.00354652f
c7 13 VSS 0.0183914f
c8 14 VSS 0.00306585f
c9 15 VSS 0.00542482f
c10 16 VSS 0.00282549f
r1 33 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 11 32 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r4 31 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r6 3 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r7 27 28 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r8 25 28 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r9 13 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r10 13 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r11 16 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r12 16 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r13 22 23 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1640 $X2=0.4590 $Y2=0.2160
r14 22 21 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1640 $X2=0.4590 $Y2=0.0920
r15 14 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r16 14 21 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0920
r17 19 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4455 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r18 15 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r19 2 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r20 10 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r21 18 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r22 1 11 1e-05
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0327274f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0425409f
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%NET041 VSS 2 3 1
c1 1 VSS 0.00100372f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3240 $Y2=0.2025
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%NET43 VSS 2 3 1
c1 1 VSS 0.000962293f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%NET015 VSS 11 17 18 2 1 8 9 7
c1 1 VSS 0.00770242f
c2 2 VSS 0.00711241f
c3 7 VSS 0.00371304f
c4 8 VSS 0.00339014f
c5 9 VSS 0.0111622f
r1 18 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 2 16 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r4 17 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r5 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r6 13 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r7 12 13 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3195
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r8 9 12 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r9 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r10 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r11 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r12 1 7 1e-05
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%B VSS 20 3 4 1 5
c1 1 VSS 0.010321f
c2 3 VSS 0.0363952f
c3 4 VSS 0.0469834f
c4 5 VSS 0.00512041f
r1 4 17 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r2 20 19 7.92845 $w=1.3e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1010
r3 5 19 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0725 $X2=0.1350 $Y2=0.1010
r4 15 17 10.5547 $w=1.466e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r5 14 15 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2845 $Y2=0.1350
r6 13 14 96.7394 $w=9.3e-09 $l=4.15e-08 $layer=LIG $thickness=4.8e-08 $X=0.2285
+ $Y=0.1350 $X2=0.2700 $Y2=0.1350
r7 12 13 97.9049 $w=9.3e-09 $l=4.2e-08 $layer=LIG $thickness=4.8e-08 $X=0.1865
+ $Y=0.1350 $X2=0.2285 $Y2=0.1350
r8 11 12 57.1112 $w=9.3e-09 $l=2.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.1620
+ $Y=0.1350 $X2=0.1865 $Y2=0.1350
r9 10 11 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.1475
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r10 8 10 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1445 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r11 7 8 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r12 20 7 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r13 1 7 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r14 1 9 1.40189 $w=1.265e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1245 $Y2=0.1350
r15 3 7 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r16 3 9 1.4802 $w=2.16633e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1245 $Y2=0.1350
r17 3 10 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%A VSS 19 5 6 1 8 14 7 10 2 11 15
c1 1 VSS 0.00463939f
c2 2 VSS 0.00410199f
c3 5 VSS 0.0713896f
c4 6 VSS 0.082565f
c5 7 VSS 0.013605f
c6 8 VSS 0.0130283f
c7 9 VSS 0.000377565f
c8 10 VSS 0.00501313f
c9 11 VSS 0.0043531f
c10 12 VSS 0.00501228f
c11 13 VSS 0.00241984f
c12 14 VSS 0.000476169f
c13 15 VSS 0.000896465f
r1 2 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r2 6 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 30 31 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1235 $X2=0.3510 $Y2=0.1350
r4 11 15 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1010 $X2=0.3510 $Y2=0.0720
r5 11 30 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1010 $X2=0.3510 $Y2=0.1235
r6 15 29 9.89378 $w=1.39091e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.3015 $Y2=0.0720
r7 10 14 4.55457 $w=1.3814e-08 $l=2.75545e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.0720 $X2=0.2160 $Y2=0.0665
r8 10 29 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0720 $X2=0.3015 $Y2=0.0720
r9 9 13 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0360
r10 9 14 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0665
r11 13 26 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1935 $Y2=0.0360
r12 25 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1935 $Y2=0.0360
r13 24 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1710 $Y2=0.0360
r14 23 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1530 $Y2=0.0360
r15 22 23 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1100
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r16 8 12 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0920 $Y=0.0360 $X2=0.0810 $Y2=0.0360
r17 8 22 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0920
+ $Y=0.0360 $X2=0.1100 $Y2=0.0360
r18 12 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0810 $Y=0.0360 $X2=0.0810 $Y2=0.0575
r19 19 7 8.62802 $w=1.3e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.0980
r20 7 21 9.44419 $w=1.3e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0980 $X2=0.0810 $Y2=0.0575
r21 5 1 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r22 19 1 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_XNOR2xp5_ASAP7_75t_R%NET29 VSS 9 34 41 42 13 4 11 12 3 1 15 16 10 17
+ 19
c1 1 VSS 0.00188329f
c2 3 VSS 0.00910568f
c3 4 VSS 0.00620993f
c4 9 VSS 0.0421538f
c5 10 VSS 0.00521645f
c6 11 VSS 0.00624721f
c7 12 VSS 0.00825779f
c8 13 VSS 0.00208184f
c9 14 VSS 0.000825941f
c10 15 VSS 0.00721881f
c11 16 VSS 0.00180817f
c12 17 VSS 0.000499583f
c13 18 VSS 0.00269255f
c14 19 VSS 0.000441598f
r1 42 40 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 3 40 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 11 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 41 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 3 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1080 $Y2=0.2340
r6 37 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r7 35 38 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r8 12 18 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1710 $Y2=0.2340
r9 12 35 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1350 $Y2=0.2340
r10 10 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r11 34 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r12 4 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1745 $Y=0.0675
+ $X2=0.1710 $Y2=0.0900
r13 14 29 2.45586 $w=1.44e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.2160 $X2=0.1710 $Y2=0.2035
r14 14 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.2160 $X2=0.1710 $Y2=0.2340
r15 30 31 9.67738 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0900 $X2=0.1710 $Y2=0.1315
r16 13 17 3.47612 $w=1.45278e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.1765 $X2=0.1710 $Y2=0.1945
r17 13 31 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1765 $X2=0.1710 $Y2=0.1315
r18 17 29 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1945 $X2=0.1710 $Y2=0.2035
r19 28 29 3.50522 $w=1.40294e-08 $l=2.31625e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1935 $Y=0.1980 $X2=0.1710 $Y2=0.2035
r20 27 28 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1980 $X2=0.1935 $Y2=0.1980
r21 26 27 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2990
+ $Y=0.1980 $X2=0.2315 $Y2=0.1980
r22 25 26 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.2990 $Y2=0.1980
r23 24 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3735
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r24 15 19 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3915 $Y=0.1980 $X2=0.4050 $Y2=0.1980
r25 15 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1980 $X2=0.3735 $Y2=0.1980
r26 19 23 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1765
r27 22 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1540 $X2=0.4050 $Y2=0.1765
r28 21 22 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1540
r29 16 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1235 $X2=0.4050 $Y2=0.1350
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r31 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends


*
.SUBCKT XNOR2xp5_ASAP7_75t_R VSS VDD A B Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* Y Y
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM5_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "XNOR2xp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "XNOR2xp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_15
cc_1 N_noxref_15_1 N_B_1 0.00113262f
cc_2 N_noxref_15_1 N_MM5_g 0.00235474f
cc_3 N_noxref_15_1 N_Y_11 0.0364567f
cc_4 N_noxref_15_1 N_noxref_13_1 0.00749686f
cc_5 N_noxref_15_1 N_noxref_14_1 0.00089527f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_12
cc_6 N_noxref_12_1 N_B_1 0.000989492f
cc_7 N_noxref_12_1 N_MM2_g 0.00227875f
cc_8 N_noxref_12_1 N_NET29_4 0.0015781f
cc_9 N_noxref_12_1 N_NET29_10 0.0368249f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_13
cc_10 N_noxref_13_1 N_B_1 0.00138309f
cc_11 N_noxref_13_1 N_MM2_g 0.00430793f
cc_12 N_noxref_13_1 N_NET29_11 0.000529488f
cc_13 N_noxref_13_1 N_noxref_12_1 0.000966724f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_14
cc_14 N_noxref_14_1 N_B_1 0.00107878f
cc_15 N_noxref_14_1 N_MM5_g 0.00230298f
cc_16 N_noxref_14_1 N_NET29_4 0.00100452f
cc_17 N_noxref_14_1 N_NET015_7 0.0351653f
cc_18 N_noxref_14_1 N_noxref_12_1 0.00731503f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_16
cc_19 N_noxref_16_1 N_MM6_g 0.00145605f
cc_20 N_noxref_16_1 N_Y_10 0.0382527f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_17
cc_21 N_noxref_17_1 N_MM6_g 0.00145686f
cc_22 N_noxref_17_1 N_Y_12 0.038395f
cc_23 N_noxref_17_1 N_noxref_16_1 0.00177384f
x_PM_XNOR2xp5_ASAP7_75t_R%Y VSS Y N_MM6_d N_MM9_d N_MM10_d N_Y_1 N_Y_11 N_Y_12
+ N_Y_3 N_Y_2 N_Y_13 N_Y_10 N_Y_14 N_Y_15 PM_XNOR2xp5_ASAP7_75t_R%Y
cc_24 N_Y_1 N_MM5_g 0.00189176f
cc_25 N_Y_11 N_B_1 0.00235336f
cc_26 N_Y_11 N_MM5_g 0.0358766f
cc_27 N_Y_12 N_MM6_g 0.0158116f
cc_28 N_Y_3 N_NET29_1 0.000893349f
cc_29 N_Y_2 N_MM6_g 0.00106929f
cc_30 N_Y_1 N_NET29_15 0.00120173f
cc_31 N_Y_3 N_MM6_g 0.00139796f
cc_32 N_Y_13 N_NET29_19 0.00163679f
cc_33 N_Y_10 N_NET29_1 0.00164114f
cc_34 N_Y_14 N_NET29_16 0.00447443f
cc_35 N_Y_13 N_NET29_15 0.0136927f
cc_36 N_Y_10 N_MM6_g 0.0546044f
cc_37 N_Y_15 N_NET015_9 0.000794603f
cc_38 N_Y_2 N_NET015_2 0.00519223f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_11
cc_39 N_noxref_11_1 N_MM3_g 0.00376903f
cc_40 N_noxref_11_1 N_noxref_10_1 0.00192672f
x_PM_XNOR2xp5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_XNOR2xp5_ASAP7_75t_R%noxref_10
cc_41 N_noxref_10_1 N_MM3_g 0.00189795f
x_PM_XNOR2xp5_ASAP7_75t_R%NET041 VSS N_MM10_s N_MM11_d N_NET041_1
+ PM_XNOR2xp5_ASAP7_75t_R%NET041
cc_42 N_NET041_1 N_MM4_g 0.0172274f
cc_43 N_NET041_1 N_MM5_g 0.0174153f
x_PM_XNOR2xp5_ASAP7_75t_R%NET43 VSS N_MM3_d N_MM2_s N_NET43_1
+ PM_XNOR2xp5_ASAP7_75t_R%NET43
cc_44 N_NET43_1 N_MM3_g 0.0172926f
cc_45 N_NET43_1 N_MM2_g 0.0172481f
x_PM_XNOR2xp5_ASAP7_75t_R%NET015 VSS N_MM5_d N_MM4_d N_MM6_s N_NET015_2
+ N_NET015_1 N_NET015_8 N_NET015_9 N_NET015_7 PM_XNOR2xp5_ASAP7_75t_R%NET015
cc_46 N_NET015_2 N_A_11 0.000617549f
cc_47 N_NET015_1 N_A_10 0.0016924f
cc_48 N_NET015_8 N_A_2 0.00077967f
cc_49 N_NET015_2 N_MM4_g 0.00129612f
cc_50 N_NET015_9 N_A_15 0.00131106f
cc_51 N_NET015_9 N_A_10 0.00800511f
cc_52 N_NET015_8 N_MM4_g 0.0344612f
cc_53 N_NET015_1 N_MM5_g 0.0015475f
cc_54 N_NET015_7 N_B_1 0.00211644f
cc_55 N_NET015_7 N_MM5_g 0.0340322f
cc_56 N_NET015_8 N_NET29_4 0.000420978f
cc_57 N_NET015_7 N_NET29_4 0.000569672f
cc_58 N_NET015_8 N_NET29_1 0.000653019f
cc_59 N_NET015_2 N_MM6_g 0.000899813f
cc_60 N_NET015_8 N_MM6_g 0.0341313f
x_PM_XNOR2xp5_ASAP7_75t_R%B VSS B N_MM2_g N_MM5_g N_B_1 N_B_5
+ PM_XNOR2xp5_ASAP7_75t_R%B
cc_61 N_B_1 N_MM3_g 0.00109758f
cc_62 N_B_1 N_A_1 0.00198128f
cc_63 N_B_5 N_A_8 0.00102986f
cc_64 N_B_1 N_A_14 0.00191491f
cc_65 N_MM5_g N_MM4_g 0.00491394f
cc_66 N_B_5 N_A_7 0.00641124f
cc_67 N_MM2_g N_MM3_g 0.00760308f
x_PM_XNOR2xp5_ASAP7_75t_R%A VSS A N_MM3_g N_MM4_g N_A_1 N_A_8 N_A_14 N_A_7
+ N_A_10 N_A_2 N_A_11 N_A_15 PM_XNOR2xp5_ASAP7_75t_R%A
x_PM_XNOR2xp5_ASAP7_75t_R%NET29 VSS N_MM6_g N_MM2_d N_MM0_d N_MM1_d N_NET29_13
+ N_NET29_4 N_NET29_11 N_NET29_12 N_NET29_3 N_NET29_1 N_NET29_15 N_NET29_16
+ N_NET29_10 N_NET29_17 N_NET29_19 PM_XNOR2xp5_ASAP7_75t_R%NET29
cc_68 N_NET29_13 N_MM3_g 0.000297871f
cc_69 N_NET29_4 N_MM3_g 0.000302229f
cc_70 N_NET29_11 N_A_1 0.00032756f
cc_71 N_NET29_12 N_A_7 0.000576303f
cc_72 N_NET29_3 N_MM3_g 0.000746496f
cc_73 N_NET29_4 N_A_10 0.000801045f
cc_74 N_NET29_1 N_A_2 0.00187579f
cc_75 N_NET29_13 N_A_7 0.00134378f
cc_76 N_NET29_13 N_A_8 0.00168739f
cc_77 N_NET29_4 N_A_8 0.00172667f
cc_78 N_NET29_15 N_A_11 0.0020469f
cc_79 N_NET29_13 N_A_14 0.00263235f
cc_80 N_MM6_g N_MM4_g 0.0033796f
cc_81 N_NET29_16 N_A_11 0.00366486f
cc_82 N_NET29_11 N_MM3_g 0.0262115f
cc_83 N_NET29_10 N_B_5 0.000297179f
cc_84 N_NET29_4 N_B_5 0.000510941f
cc_85 N_NET29_17 N_B_5 0.000703189f
cc_86 N_NET29_13 N_B_1 0.000705954f
cc_87 N_NET29_3 N_MM2_g 0.000706997f
cc_88 N_NET29_12 N_B_5 0.000827021f
cc_89 N_NET29_15 N_B_1 0.000890937f
cc_90 N_NET29_4 N_MM2_g 0.00310587f
cc_91 N_NET29_11 N_MM2_g 0.0109859f
cc_92 N_NET29_4 N_B_1 0.00485262f
cc_93 N_NET29_13 N_B_5 0.0113616f
cc_94 N_NET29_10 N_MM2_g 0.0501545f
*END of XNOR2xp5_ASAP7_75t_R.pxi
.ENDS
** Design:	MAJIxp5_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "MAJIxp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "MAJIxp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_MAJIxp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.0425213f
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%NET17 VSS 2 3 1
c1 1 VSS 0.00100423f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2160 $Y2=0.0675
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.042448f
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000985874f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2160 $Y2=0.2025
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%C VSS 17 3 4 5 1
c1 1 VSS 0.0155361f
c2 3 VSS 0.0826232f
c3 4 VSS 0.086442f
c4 5 VSS 0.00483065f
r1 4 14 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 17 18 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1160 $X2=0.1350 $Y2=0.1212
r3 5 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r4 5 18 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1212
r5 12 14 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1765 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 11 12 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1765 $Y2=0.1350
r7 10 11 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r8 8 10 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.1445
+ $Y=0.1350 $X2=0.1475 $Y2=0.1350
r9 7 8 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r10 1 7 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r11 1 9 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1245 $Y2=0.1350
r12 3 7 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r13 3 9 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1 $thickness=5.5619e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1245 $Y2=0.1350
r14 3 10 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%B VSS 18 5 6 12 1 9 2 11 15 10 7 16
c1 1 VSS 0.00425445f
c2 2 VSS 0.000492087f
c3 5 VSS 0.0804219f
c4 6 VSS 0.00634214f
c5 7 VSS 0.0156656f
c6 8 VSS 0.00576573f
c7 9 VSS 0.00353914f
c8 10 VSS 0.00888536f
c9 11 VSS 0.00200068f
c10 12 VSS 0.00247873f
c11 13 VSS 0.00295784f
c12 14 VSS 0.00457223f
c13 15 VSS 0.00102152f
c14 16 VSS 0.000626249f
r1 2 32 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r2 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r3 12 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r4 12 15 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2160 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 15 31 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1540
r6 11 16 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1765 $X2=0.1890 $Y2=0.1980
r7 11 31 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1540
r8 16 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1980 $X2=0.1620 $Y2=0.1980
r9 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1980 $X2=0.1620 $Y2=0.1980
r10 28 29 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1105
+ $Y=0.1980 $X2=0.1350 $Y2=0.1980
r11 27 28 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.1980 $X2=0.1105 $Y2=0.1980
r12 10 14 7.2121 $w=1.41842e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0650 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r13 10 27 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.0650
+ $Y=0.1980 $X2=0.0945 $Y2=0.1980
r14 14 26 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r15 8 13 3.2503 $w=1.53684e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1540 $X2=0.0270 $Y2=0.1350
r16 8 26 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1540 $X2=0.0270 $Y2=0.1765
r17 7 13 7.44771 $w=1.42162e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0980 $X2=0.0270 $Y2=0.1350
r18 19 20 3.08976 $w=1.3e-08 $l=1.33e-08 $layer=M1 $thickness=3.6e-08 $X=0.0677
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r19 18 19 1.10765 $w=1.3e-08 $l=4.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.0630
+ $Y=0.1350 $X2=0.0677 $Y2=0.1350
r20 18 9 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.0630
+ $Y=0.1350 $X2=0.0492 $Y2=0.1350
r21 9 13 4.00816 $w=1.50225e-08 $l=2.22e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0492 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r22 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r23 1 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%NET1 VSS 12 13 24 7 1 9 8 2
c1 1 VSS 0.010186f
c2 2 VSS 0.00542391f
c3 7 VSS 0.00471491f
c4 8 VSS 0.00264525f
c5 9 VSS 0.0258804f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.0675 $X2=0.3220 $Y2=0.0675
r2 24 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.0675 $X2=0.3095 $Y2=0.0675
r3 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.0675
+ $X2=0.3240 $Y2=0.0360
r4 20 21 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2850
+ $Y=0.0360 $X2=0.3240 $Y2=0.0360
r5 19 20 15.7403 $w=1.3e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.2175
+ $Y=0.0360 $X2=0.2850 $Y2=0.0360
r6 18 19 12.942 $w=1.3e-08 $l=5.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2175 $Y2=0.0360
r7 17 18 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r8 16 17 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1215
+ $Y=0.0360 $X2=0.1350 $Y2=0.0360
r9 15 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r10 14 15 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0970
+ $Y=0.0360 $X2=0.1080 $Y2=0.0360
r11 9 14 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0945
+ $Y=0.0360 $X2=0.0970 $Y2=0.0360
r12 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r13 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r14 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r15 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r16 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00569877f
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00590537f
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%Y VSS 25 16 17 36 37 9 2 1 8 10 7 11 12 13
c1 1 VSS 0.00364802f
c2 2 VSS 0.00358233f
c3 7 VSS 0.00301191f
c4 8 VSS 0.00269556f
c5 9 VSS 0.000925435f
c6 10 VSS 0.000793611f
c7 11 VSS 0.00126635f
c8 12 VSS 0.000733969f
c9 13 VSS 0.000740498f
r1 37 35 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 35 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 36 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2690 $Y2=0.1980
r6 31 32 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2690
+ $Y=0.1980 $X2=0.2830 $Y2=0.1980
r7 29 32 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1980 $X2=0.2830 $Y2=0.1980
r8 28 29 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.1980 $X2=0.2970 $Y2=0.1980
r9 10 13 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3405 $Y=0.1980 $X2=0.3520 $Y2=0.1980
r10 10 28 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3405
+ $Y=0.1980 $X2=0.3220 $Y2=0.1980
r11 13 27 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3520 $Y=0.1980 $X2=0.3520 $Y2=0.1765
r12 26 27 6.70421 $w=1.3e-08 $l=2.88e-08 $layer=M1 $thickness=3.6e-08 $X=0.3520
+ $Y=0.1477 $X2=0.3520 $Y2=0.1765
r13 25 26 3.90593 $w=1.3e-08 $l=1.67e-08 $layer=M1 $thickness=3.6e-08 $X=0.3520
+ $Y=0.1310 $X2=0.3520 $Y2=0.1477
r14 25 24 2.97317 $w=1.3e-08 $l=1.28e-08 $layer=M1 $thickness=3.6e-08 $X=0.3520
+ $Y=0.1310 $X2=0.3520 $Y2=0.1182
r15 11 12 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3520 $Y=0.0935 $X2=0.3520 $Y2=0.0720
r16 11 24 5.77145 $w=1.3e-08 $l=2.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.3520
+ $Y=0.0935 $X2=0.3520 $Y2=0.1182
r17 12 23 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3520 $Y=0.0720 $X2=0.3405 $Y2=0.0720
r18 22 23 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.3220
+ $Y=0.0720 $X2=0.3405 $Y2=0.0720
r19 21 22 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.0720 $X2=0.3220 $Y2=0.0720
r20 20 21 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2830
+ $Y=0.0720 $X2=0.2970 $Y2=0.0720
r21 19 20 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2690
+ $Y=0.0720 $X2=0.2830 $Y2=0.0720
r22 18 19 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0720 $X2=0.2690 $Y2=0.0720
r23 9 18 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2560
+ $Y=0.0720 $X2=0.2585 $Y2=0.0720
r24 1 19 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2690 $Y2=0.0720
r25 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r26 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r27 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r28 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%NET3 VSS 12 13 21 7 1 9 8 2
c1 1 VSS 0.0100554f
c2 2 VSS 0.00536451f
c3 7 VSS 0.00463203f
c4 8 VSS 0.00261844f
c5 9 VSS 0.0221353f
r1 8 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3095 $Y=0.2025 $X2=0.3220 $Y2=0.2025
r2 21 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3095 $Y2=0.2025
r3 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3240 $Y=0.2025
+ $X2=0.3240 $Y2=0.2340
r4 17 18 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2850
+ $Y=0.2340 $X2=0.3240 $Y2=0.2340
r5 16 17 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2265
+ $Y=0.2340 $X2=0.2850 $Y2=0.2340
r6 15 16 16.0901 $w=1.3e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1575
+ $Y=0.2340 $X2=0.2265 $Y2=0.2340
r7 14 15 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1575 $Y2=0.2340
r8 9 14 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0965
+ $Y=0.2340 $X2=0.1080 $Y2=0.2340
r9 1 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r10 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r11 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r12 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r13 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
.ends

.subckt PM_MAJIxp5_ASAP7_75t_R%A VSS 7 3 1 4
c1 1 VSS 0.00900255f
c2 3 VSS 0.00890853f
c3 4 VSS 0.00487235f
r1 7 8 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1160 $X2=0.2970 $Y2=0.1212
r2 4 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1212
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends


*
.SUBCKT MAJIxp5_ASAP7_75t_R VSS VDD B C A Y
*
* VSS VSS
* VDD VDD
* B B
* C C
* A A
* Y Y
*
*

MM1 N_MM1_d N_MM1_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM0_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "MAJIxp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "MAJIxp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_MAJIxp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_MAJIxp5_ASAP7_75t_R%noxref_12
cc_1 N_noxref_12_1 N_MM1_g 0.00217576f
cc_2 N_noxref_12_1 N_noxref_11_1 0.00177466f
x_PM_MAJIxp5_ASAP7_75t_R%NET17 VSS N_MM4_d N_MM3_s N_NET17_1
+ PM_MAJIxp5_ASAP7_75t_R%NET17
cc_3 N_NET17_1 N_MM3_g 0.0172525f
cc_4 N_NET17_1 N_MM4_g 0.0174726f
x_PM_MAJIxp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_MAJIxp5_ASAP7_75t_R%noxref_11
cc_5 N_noxref_11_1 N_MM1_g 0.00221502f
x_PM_MAJIxp5_ASAP7_75t_R%NET16 VSS N_MM9_d N_MM8_s N_NET16_1
+ PM_MAJIxp5_ASAP7_75t_R%NET16
cc_6 N_NET16_1 N_MM3_g 0.0172156f
cc_7 N_NET16_1 N_MM4_g 0.0173778f
x_PM_MAJIxp5_ASAP7_75t_R%C VSS C N_MM2_g N_MM4_g N_C_5 N_C_1
+ PM_MAJIxp5_ASAP7_75t_R%C
cc_8 N_MM4_g N_B_12 0.000449542f
cc_9 N_MM4_g N_B_1 0.000451453f
cc_10 N_MM4_g N_B_9 0.000636201f
cc_11 N_MM4_g N_B_2 0.000639569f
cc_12 N_C_5 N_B_11 0.000803694f
cc_13 N_C_5 N_B_15 0.000822224f
cc_14 N_C_5 N_B_10 0.00132851f
cc_15 N_C_1 N_B_15 0.00222023f
cc_16 N_MM2_g N_MM1_g 0.00338752f
cc_17 N_C_5 N_B_9 0.00446017f
cc_18 N_MM4_g N_MM3_g 0.00764704f
x_PM_MAJIxp5_ASAP7_75t_R%B VSS B N_MM1_g N_MM3_g N_B_12 N_B_1 N_B_9 N_B_2
+ N_B_11 N_B_15 N_B_10 N_B_7 N_B_16 PM_MAJIxp5_ASAP7_75t_R%B
x_PM_MAJIxp5_ASAP7_75t_R%NET1 VSS N_MM1_d N_MM2_d N_MM0_s N_NET1_7 N_NET1_1
+ N_NET1_9 N_NET1_8 N_NET1_2 PM_MAJIxp5_ASAP7_75t_R%NET1
cc_19 N_NET1_7 N_B_7 0.000434857f
cc_20 N_NET1_7 N_B_1 0.00068017f
cc_21 N_NET1_1 N_MM1_g 0.00104965f
cc_22 N_NET1_9 N_B_12 0.00122558f
cc_23 N_NET1_7 N_MM1_g 0.0350445f
cc_24 N_NET1_1 N_MM2_g 0.00126885f
cc_25 N_NET1_9 N_C_5 0.00144076f
cc_26 N_NET1_1 N_C_5 0.00189058f
cc_27 N_NET1_7 N_MM2_g 0.0352624f
cc_28 N_NET1_8 N_A_1 0.000722956f
cc_29 N_NET1_2 N_MM0_g 0.00102492f
cc_30 N_NET1_8 N_MM0_g 0.0344853f
x_PM_MAJIxp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_MAJIxp5_ASAP7_75t_R%noxref_13
cc_31 N_noxref_13_1 N_MM0_g 0.00144423f
cc_32 N_noxref_13_1 N_NET1_8 0.0363826f
cc_33 N_noxref_13_1 N_NET3_8 0.000472185f
cc_34 N_noxref_13_1 N_Y_7 0.000726864f
x_PM_MAJIxp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_MAJIxp5_ASAP7_75t_R%noxref_14
cc_35 N_noxref_14_1 N_MM0_g 0.00143979f
cc_36 N_noxref_14_1 N_NET1_8 0.000476144f
cc_37 N_noxref_14_1 N_NET3_8 0.0361761f
cc_38 N_noxref_14_1 N_Y_8 0.000727239f
cc_39 N_noxref_14_1 N_noxref_13_1 0.00177174f
x_PM_MAJIxp5_ASAP7_75t_R%Y VSS Y N_MM3_d N_MM0_d N_MM8_d N_MM5_d N_Y_9 N_Y_2
+ N_Y_1 N_Y_8 N_Y_10 N_Y_7 N_Y_11 N_Y_12 N_Y_13 PM_MAJIxp5_ASAP7_75t_R%Y
cc_40 N_Y_9 N_B_12 0.00049802f
cc_41 N_Y_2 N_B_2 0.000768448f
cc_42 N_Y_1 N_MM3_g 0.00118327f
cc_43 N_Y_2 N_MM3_g 0.00125039f
cc_44 N_Y_8 N_B_2 0.00161739f
cc_45 N_Y_10 N_B_12 0.00168971f
cc_46 N_Y_8 N_MM3_g 0.0151144f
cc_47 N_Y_7 N_MM3_g 0.054754f
cc_48 N_Y_2 N_A_1 0.000837342f
cc_49 N_Y_1 N_MM0_g 0.000888968f
cc_50 N_Y_2 N_MM0_g 0.000889984f
cc_51 N_Y_10 N_A_4 0.00110857f
cc_52 N_Y_9 N_A_4 0.00115507f
cc_53 N_Y_8 N_A_1 0.00155895f
cc_54 N_Y_11 N_A_4 0.00456306f
cc_55 N_Y_8 N_MM0_g 0.0148926f
cc_56 N_Y_7 N_MM0_g 0.0528616f
cc_57 N_Y_12 N_NET1_9 0.0006069f
cc_58 N_Y_9 N_NET1_2 0.000644131f
cc_59 N_Y_7 N_NET1_8 0.000679579f
cc_60 N_Y_11 N_NET1_2 0.000684527f
cc_61 N_Y_1 N_NET1_2 0.00418149f
cc_62 N_Y_9 N_NET1_9 0.00944163f
cc_63 N_Y_13 N_NET3_9 0.000605682f
cc_64 N_Y_10 N_NET3_2 0.00064116f
cc_65 N_Y_11 N_NET3_2 0.000658939f
cc_66 N_Y_8 N_NET3_8 0.000680046f
cc_67 N_Y_2 N_NET3_2 0.00414893f
cc_68 N_Y_10 N_NET3_9 0.00914447f
x_PM_MAJIxp5_ASAP7_75t_R%NET3 VSS N_MM6_d N_MM7_d N_MM5_s N_NET3_7 N_NET3_1
+ N_NET3_9 N_NET3_8 N_NET3_2 PM_MAJIxp5_ASAP7_75t_R%NET3
cc_69 N_NET3_7 N_B_10 0.000398974f
cc_70 N_NET3_7 N_B_1 0.000691871f
cc_71 N_NET3_1 N_MM1_g 0.00163445f
cc_72 N_NET3_9 N_B_10 0.00442606f
cc_73 N_NET3_9 N_B_16 0.0053591f
cc_74 N_NET3_7 N_MM1_g 0.0347295f
cc_75 N_NET3_1 N_MM2_g 0.000929125f
cc_76 N_NET3_7 N_MM2_g 0.0351857f
cc_77 N_NET3_8 N_A_1 0.00076267f
cc_78 N_NET3_2 N_MM0_g 0.00101062f
cc_79 N_NET3_8 N_MM0_g 0.0342473f
x_PM_MAJIxp5_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_MAJIxp5_ASAP7_75t_R%A
cc_80 N_A_1 N_B_2 0.000886983f
cc_81 N_A_4 N_B_12 0.00169977f
cc_82 N_MM0_g N_MM3_g 0.00413988f
*END of MAJIxp5_ASAP7_75t_R.pxi
.ENDS
** Design:	MAJx2_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "MAJx2_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "MAJx2_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_MAJx2_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.0423307f
.ends

.subckt PM_MAJx2_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.0423307f
.ends

.subckt PM_MAJx2_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00571289f
.ends

.subckt PM_MAJx2_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00584057f
.ends

.subckt PM_MAJx2_ASAP7_75t_R%NET17 VSS 2 3 1
c1 1 VSS 0.00099779f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_MAJx2_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.00100152f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_MAJx2_ASAP7_75t_R%Y VSS 22 16 17 32 33 10 7 8 9 11 1 2
c1 1 VSS 0.010194f
c2 2 VSS 0.0105571f
c3 7 VSS 0.00450404f
c4 8 VSS 0.00450982f
c5 9 VSS 0.00898504f
c6 10 VSS 0.00936981f
c7 11 VSS 0.00734686f
c8 12 VSS 0.00349051f
c9 13 VSS 0.00355402f
r1 33 31 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r2 2 31 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r4 32 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r5 2 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3775 $Y2=0.2340
r6 10 26 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r7 10 28 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.2340 $X2=0.3775 $Y2=0.2340
r8 13 25 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r9 13 26 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4185 $Y2=0.2340
r10 24 25 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4590 $Y2=0.2160
r11 23 24 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1485 $X2=0.4590 $Y2=0.1780
r12 22 23 0.23319 $w=1.3e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1485
r13 22 21 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1050
r14 11 12 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r15 11 21 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.1050
r16 12 20 7.79507 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4185 $Y2=0.0360
r17 19 20 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r18 18 19 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3775
+ $Y=0.0360 $X2=0.3865 $Y2=0.0360
r19 9 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.0360 $X2=0.3775 $Y2=0.0360
r20 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3775 $Y2=0.0360
r21 17 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r22 1 15 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r23 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r24 16 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
.ends

.subckt PM_MAJx2_ASAP7_75t_R%C VSS 17 3 4 5 1
c1 1 VSS 0.0154146f
c2 3 VSS 0.0854816f
c3 4 VSS 0.0826398f
c4 5 VSS 0.00362955f
r1 3 13 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r2 17 18 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1212
r3 5 7 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r4 5 18 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1212
r5 11 13 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2015 $Y=0.1350 $X2=0.1890 $Y2=0.1350
r6 10 11 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2160 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r7 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2305
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r8 8 15 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.2525
+ $Y=0.1350 $X2=0.2535 $Y2=0.1350
r9 7 8 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2525 $Y2=0.1350
r10 1 7 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r11 1 9 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2305 $Y2=0.1350
r12 4 7 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r13 4 9 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.2430 $Y=0.1350 $X2=0.2305 $Y2=0.1350
r14 4 15 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.2430 $Y=0.1350 $X2=0.2535 $Y2=0.1350
.ends

.subckt PM_MAJx2_ASAP7_75t_R%NET1 VSS 11 18 19 7 1 8 2 9
c1 1 VSS 0.00531144f
c2 2 VSS 0.0100647f
c3 7 VSS 0.00262752f
c4 8 VSS 0.00459542f
c5 9 VSS 0.0226021f
r1 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 2 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r4 18 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r5 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r6 13 14 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r7 12 13 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r8 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r9 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r10 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r11 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r12 1 7 1e-05
.ends

.subckt PM_MAJx2_ASAP7_75t_R%MAJI VSS 9 10 50 51 62 63 12 3 4 15 14 13 11 1 16
+ 17 18 19
c1 1 VSS 0.00725807f
c2 3 VSS 0.0034703f
c3 4 VSS 0.00354572f
c4 9 VSS 0.0805051f
c5 10 VSS 0.0808278f
c6 11 VSS 0.00459227f
c7 12 VSS 0.00463052f
c8 13 VSS 0.00419076f
c9 14 VSS 0.00940196f
c10 15 VSS 0.00140822f
c11 16 VSS 0.00194021f
c12 17 VSS 0.00162106f
c13 18 VSS 0.00161057f
c14 19 VSS 0.000480903f
r1 63 61 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 4 61 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 12 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 62 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 4 57 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1090 $Y2=0.1980
r6 56 57 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.1980 $X2=0.1090 $Y2=0.1980
r7 55 56 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0950 $Y2=0.1980
r8 54 55 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 15 18 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0380 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 15 54 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0380
+ $Y=0.1980 $X2=0.0560 $Y2=0.1980
r11 18 53 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r12 52 53 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1765
r13 13 17 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0935 $X2=0.0270 $Y2=0.0720
r14 13 52 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0935 $X2=0.0270 $Y2=0.1350
r15 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r16 3 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r17 11 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r18 50 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r19 17 47 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0720 $X2=0.0380 $Y2=0.0720
r20 3 43 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1090 $Y2=0.0720
r21 46 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.0720 $X2=0.0380 $Y2=0.0720
r22 45 46 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0560 $Y2=0.0720
r23 43 44 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1090
+ $Y=0.0720 $X2=0.1195 $Y2=0.0720
r24 42 43 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.0720 $X2=0.1090 $Y2=0.0720
r25 42 45 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.0720 $X2=0.0810 $Y2=0.0720
r26 41 44 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1595
+ $Y=0.0720 $X2=0.1195 $Y2=0.0720
r27 40 41 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.1595 $Y2=0.0720
r28 39 40 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r29 38 39 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2675
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r30 37 38 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0720 $X2=0.2675 $Y2=0.0720
r31 36 37 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2995
+ $Y=0.0720 $X2=0.2835 $Y2=0.0720
r32 35 36 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0720 $X2=0.2995 $Y2=0.0720
r33 34 35 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3485
+ $Y=0.0720 $X2=0.3240 $Y2=0.0720
r34 14 19 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3660 $Y=0.0720 $X2=0.3770 $Y2=0.0720
r35 14 34 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3660
+ $Y=0.0720 $X2=0.3485 $Y2=0.0720
r36 19 32 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3770 $Y=0.0720 $X2=0.3770 $Y2=0.0935
r37 10 28 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r38 16 30 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3770
+ $Y=0.1160 $X2=0.3770 $Y2=0.1350
r39 16 32 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3770
+ $Y=0.1160 $X2=0.3770 $Y2=0.0935
r40 26 28 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r41 25 26 2.65825 $w=1.53e-08 $l=4.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3880 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r42 24 25 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3770 $Y=0.1350 $X2=0.3880 $Y2=0.1350
r43 24 30 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3770 $Y=0.1350
+ $X2=0.3770 $Y2=0.1350
r44 23 24 5.90723 $w=1.53e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3670
+ $Y=0.1350 $X2=0.3770 $Y2=0.1350
r45 22 23 2.06753 $w=1.53e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3670 $Y2=0.1350
r46 9 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r47 1 21 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r48 1 22 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r49 9 21 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r50 9 22 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
.ends

.subckt PM_MAJx2_ASAP7_75t_R%A VSS 7 3 1 4
c1 1 VSS 0.00819683f
c2 3 VSS 0.00849325f
c3 4 VSS 0.00443528f
r1 7 8 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1212
r2 4 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1212
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r4 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_MAJx2_ASAP7_75t_R%NET3 VSS 12 13 21 7 1 2 8 9
c1 1 VSS 0.00543334f
c2 2 VSS 0.00997719f
c3 7 VSS 0.00262245f
c4 8 VSS 0.00462025f
c5 9 VSS 0.0243537f
r1 21 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 7 20 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 18 19 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0930 $Y2=0.2340
r5 16 19 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1515
+ $Y=0.2340 $X2=0.0930 $Y2=0.2340
r6 9 14 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2205
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r7 9 16 16.0901 $w=1.3e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2205
+ $Y=0.2340 $X2=0.1515 $Y2=0.2340
r8 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r9 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r10 2 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r11 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r12 12 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r13 1 7 1e-05
.ends

.subckt PM_MAJx2_ASAP7_75t_R%B VSS 22 5 6 7 13 11 1 8 9 10 2 14 12 15
c1 1 VSS 0.00339099f
c2 2 VSS 0.00690085f
c3 5 VSS 0.00786879f
c4 6 VSS 0.0816057f
c5 7 VSS 0.00203959f
c6 8 VSS 0.00230929f
c7 9 VSS 0.00463705f
c8 10 VSS 0.00265132f
c9 11 VSS 0.00178266f
c10 12 VSS 0.00208376f
c11 13 VSS 0.0018928f
c12 14 VSS 0.00219075f
c13 15 VSS 0.00272768f
r1 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r4 7 29 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1245
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 11 28 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1540
r6 11 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r7 8 12 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1765 $X2=0.1890 $Y2=0.1980
r8 8 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1540
r9 12 27 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1980 $X2=0.2160 $Y2=0.1980
r10 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r11 25 26 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2675
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r12 24 25 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.1980 $X2=0.2675 $Y2=0.1980
r13 22 23 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.2890
+ $Y=0.1980 $X2=0.3022 $Y2=0.1980
r14 22 9 0.641272 $w=1.3e-08 $l=2.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2890
+ $Y=0.1980 $X2=0.2862 $Y2=0.1980
r15 9 24 0.641272 $w=1.3e-08 $l=2.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2862
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r16 15 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.3240 $Y2=0.1765
r17 15 23 3.42276 $w=1.5069e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.3022 $Y2=0.1980
r18 20 21 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1565 $X2=0.3240 $Y2=0.1765
r19 10 14 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1465 $X2=0.3240 $Y2=0.1350
r20 10 20 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1465 $X2=0.3240 $Y2=0.1565
r21 14 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3105 $Y2=0.1350
r22 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3105 $Y2=0.1350
r23 13 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r24 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r25 2 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends


*
.SUBCKT MAJx2_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM11@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM0_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "MAJx2_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "MAJx2_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_MAJx2_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_MAJx2_ASAP7_75t_R%noxref_14
cc_1 N_noxref_14_1 N_MM11@2_g 0.00146601f
cc_2 N_noxref_14_1 N_Y_7 0.000843342f
x_PM_MAJx2_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_MAJx2_ASAP7_75t_R%noxref_15
cc_3 N_noxref_15_1 N_MM11@2_g 0.00147188f
cc_4 N_noxref_15_1 N_Y_8 0.000843744f
cc_5 N_noxref_15_1 N_noxref_14_1 0.00177098f
x_PM_MAJx2_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_MAJx2_ASAP7_75t_R%noxref_12
cc_6 N_noxref_12_1 N_MM0_g 0.00144364f
cc_7 N_noxref_12_1 N_MAJI_11 0.000734647f
cc_8 N_noxref_12_1 N_NET1_7 0.0363359f
cc_9 N_noxref_12_1 N_NET3_7 0.000471668f
x_PM_MAJx2_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_MAJx2_ASAP7_75t_R%noxref_13
cc_10 N_noxref_13_1 N_MM0_g 0.00145075f
cc_11 N_noxref_13_1 N_MAJI_12 0.000733669f
cc_12 N_noxref_13_1 N_NET1_7 0.000474288f
cc_13 N_noxref_13_1 N_NET3_7 0.0361995f
cc_14 N_noxref_13_1 N_noxref_12_1 0.00176881f
x_PM_MAJx2_ASAP7_75t_R%NET17 VSS N_MM3_s N_MM4_d N_NET17_1
+ PM_MAJx2_ASAP7_75t_R%NET17
cc_15 N_NET17_1 N_MM3_g 0.0172241f
cc_16 N_NET17_1 N_MM4_g 0.0174268f
x_PM_MAJx2_ASAP7_75t_R%NET16 VSS N_MM8_s N_MM9_d N_NET16_1
+ PM_MAJx2_ASAP7_75t_R%NET16
cc_17 N_NET16_1 N_MM3_g 0.0172813f
cc_18 N_NET16_1 N_MM4_g 0.0174474f
x_PM_MAJx2_ASAP7_75t_R%Y VSS Y N_MM10_d N_MM10@2_d N_MM11_d N_MM11@2_d N_Y_10
+ N_Y_7 N_Y_8 N_Y_9 N_Y_11 N_Y_1 N_Y_2 PM_MAJx2_ASAP7_75t_R%Y
cc_19 N_Y_10 N_B_15 0.00264775f
cc_20 N_Y_7 N_MAJI_1 0.000778965f
cc_21 N_Y_8 N_MM11@2_g 0.030875f
cc_22 N_Y_9 N_MAJI_14 0.00121335f
cc_23 N_Y_11 N_MAJI_1 0.00131121f
cc_24 N_Y_1 N_MAJI_16 0.00163773f
cc_25 N_Y_2 N_MM11@2_g 0.00202561f
cc_26 N_Y_1 N_MM11@2_g 0.00259591f
cc_27 N_Y_9 N_MAJI_19 0.00311176f
cc_28 N_Y_8 N_MAJI_1 0.00437087f
cc_29 N_Y_7 N_MM11_g 0.0372285f
cc_30 N_Y_7 N_MM11@2_g 0.0690284f
x_PM_MAJx2_ASAP7_75t_R%C VSS C N_MM4_g N_MM7_g N_C_5 N_C_1
+ PM_MAJx2_ASAP7_75t_R%C
cc_31 N_MM4_g N_B_13 0.000633092f
cc_32 N_C_5 N_B_11 0.000682114f
cc_33 N_C_1 N_B_1 0.000688856f
cc_34 N_C_5 N_B_8 0.000774058f
cc_35 N_C_5 N_B_9 0.00127007f
cc_36 N_C_1 N_B_11 0.00209491f
cc_37 N_MM7_g N_MM6_g 0.00337975f
cc_38 N_C_5 N_B_13 0.00355978f
cc_39 N_MM4_g N_MM3_g 0.00831749f
x_PM_MAJx2_ASAP7_75t_R%NET1 VSS N_MM0_s N_MM2_d N_MM1_d N_NET1_7 N_NET1_1
+ N_NET1_8 N_NET1_2 N_NET1_9 PM_MAJx2_ASAP7_75t_R%NET1
cc_40 N_NET1_7 N_A_1 0.000744156f
cc_41 N_NET1_1 N_MM0_g 0.0010123f
cc_42 N_NET1_7 N_MM0_g 0.0343901f
cc_43 N_NET1_8 N_B_2 0.000775684f
cc_44 N_NET1_2 N_MM6_g 0.000878668f
cc_45 N_NET1_8 N_MM6_g 0.0346991f
cc_46 N_NET1_2 N_MM7_g 0.000920115f
cc_47 N_NET1_8 N_MM7_g 0.0351918f
cc_48 N_NET1_7 N_MAJI_11 0.00126838f
cc_49 N_NET1_9 N_MAJI_17 0.000637631f
cc_50 N_NET1_1 N_MAJI_13 0.000668954f
cc_51 N_NET1_2 N_MAJI_14 0.000770027f
cc_52 N_NET1_1 N_MAJI_3 0.00412206f
cc_53 N_NET1_9 N_MAJI_14 0.0220562f
x_PM_MAJx2_ASAP7_75t_R%MAJI VSS N_MM11_g N_MM11@2_g N_MM0_d N_MM3_d N_MM5_d
+ N_MM8_d N_MAJI_12 N_MAJI_3 N_MAJI_4 N_MAJI_15 N_MAJI_14 N_MAJI_13 N_MAJI_11
+ N_MAJI_1 N_MAJI_16 N_MAJI_17 N_MAJI_18 N_MAJI_19 PM_MAJx2_ASAP7_75t_R%MAJI
cc_54 N_MAJI_12 N_MM0_g 0.0155589f
cc_55 N_MAJI_3 N_MM0_g 0.000910145f
cc_56 N_MAJI_4 N_MM0_g 0.000910195f
cc_57 N_MAJI_3 N_A_1 0.00100546f
cc_58 N_MAJI_15 N_A_4 0.00110712f
cc_59 N_MAJI_14 N_A_4 0.00121579f
cc_60 N_MAJI_12 N_A_1 0.00159919f
cc_61 N_MAJI_13 N_A_4 0.00492087f
cc_62 N_MAJI_11 N_MM0_g 0.0539369f
cc_63 N_MAJI_15 N_MM3_g 0.000213609f
cc_64 N_MAJI_4 N_MM3_g 0.00149558f
cc_65 N_MAJI_1 N_MM3_g 0.000617421f
cc_66 N_MAJI_15 N_B_8 0.000343362f
cc_67 N_MAJI_14 N_B_13 0.000457344f
cc_68 N_MAJI_12 N_MM3_g 0.0158856f
cc_69 N_MAJI_15 N_B_7 0.000617866f
cc_70 N_MAJI_16 N_B_10 0.000666347f
cc_71 N_MAJI_3 N_B_1 0.000846912f
cc_72 N_MAJI_1 N_B_2 0.00112415f
cc_73 N_MAJI_3 N_MM3_g 0.00117149f
cc_74 N_MAJI_14 N_B_14 0.00154129f
cc_75 N_MAJI_14 N_B_7 0.00164652f
cc_76 N_MAJI_16 N_B_14 0.00167899f
cc_77 N_MAJI_12 N_B_1 0.00179921f
cc_78 N_MM11_g N_MM6_g 0.00331243f
cc_79 N_MAJI_14 N_B_11 0.00365361f
cc_80 N_MAJI_11 N_MM3_g 0.0553205f
cc_81 N_MAJI_11 N_C_5 0.000517825f
cc_82 N_MAJI_14 N_C_5 0.00422198f
x_PM_MAJx2_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_MAJx2_ASAP7_75t_R%A
x_PM_MAJx2_ASAP7_75t_R%NET3 VSS N_MM7_d N_MM6_d N_MM5_s N_NET3_7 N_NET3_1
+ N_NET3_2 N_NET3_8 N_NET3_9 PM_MAJx2_ASAP7_75t_R%NET3
cc_83 N_NET3_7 N_A_1 0.000775779f
cc_84 N_NET3_1 N_MM0_g 0.00101176f
cc_85 N_NET3_7 N_MM0_g 0.0342968f
cc_86 N_NET3_2 N_B_9 0.00051712f
cc_87 N_NET3_8 N_B_2 0.000728238f
cc_88 N_NET3_2 N_MM6_g 0.00164406f
cc_89 N_NET3_9 N_B_9 0.00417248f
cc_90 N_NET3_9 N_B_12 0.0058345f
cc_91 N_NET3_8 N_MM6_g 0.0348366f
cc_92 N_NET3_2 N_MM7_g 0.000937075f
cc_93 N_NET3_8 N_MM7_g 0.0351216f
cc_94 N_NET3_9 N_MAJI_12 0.00059561f
cc_95 N_NET3_1 N_MAJI_15 0.000621844f
cc_96 N_NET3_9 N_MAJI_18 0.000639778f
cc_97 N_NET3_7 N_MAJI_12 0.000677837f
cc_98 N_NET3_1 N_MAJI_13 0.000713064f
cc_99 N_NET3_1 N_MAJI_4 0.00412823f
cc_100 N_NET3_9 N_MAJI_15 0.00874355f
x_PM_MAJx2_ASAP7_75t_R%B VSS B N_MM3_g N_MM6_g N_B_7 N_B_13 N_B_11 N_B_1 N_B_8
+ N_B_9 N_B_10 N_B_2 N_B_14 N_B_12 N_B_15 PM_MAJx2_ASAP7_75t_R%B
cc_101 N_MM3_g N_A_1 0.000847344f
cc_102 N_B_7 N_A_4 0.00172757f
cc_103 N_MM3_g N_MM0_g 0.00418692f
*END of MAJx2_ASAP7_75t_R.pxi
.ENDS
** Design:	MAJx3_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "MAJx3_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "MAJx3_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_MAJx3_ASAP7_75t_R%NET17 VSS 2 3 1
c1 1 VSS 0.000984193f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_MAJx3_ASAP7_75t_R%NET16 VSS 2 3 1
c1 1 VSS 0.000996218f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_MAJx3_ASAP7_75t_R%C VSS 18 3 4 5 1
c1 1 VSS 0.0155785f
c2 3 VSS 0.085495f
c3 4 VSS 0.0826401f
c4 5 VSS 0.00359933f
r1 18 19 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1160 $X2=0.2430 $Y2=0.1212
r2 5 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
r3 5 19 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1212
r4 4 13 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r5 12 13 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2335
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r6 10 12 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.2305 $Y=0.1350 $X2=0.2335 $Y2=0.1350
r7 9 10 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2160
+ $Y=0.1350 $X2=0.2305 $Y2=0.1350
r8 8 9 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2015
+ $Y=0.1350 $X2=0.2160 $Y2=0.1350
r9 3 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r10 1 7 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r11 1 8 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
r12 3 7 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1 $thickness=5.5619e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1785 $Y2=0.1350
r13 3 8 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1890 $Y=0.1350 $X2=0.2015 $Y2=0.1350
.ends

.subckt PM_MAJx3_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00596481f
.ends

.subckt PM_MAJx3_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00569657f
.ends

.subckt PM_MAJx3_ASAP7_75t_R%NET3 VSS 12 13 21 7 1 2 8 9
c1 1 VSS 0.00519205f
c2 2 VSS 0.0100579f
c3 7 VSS 0.00262653f
c4 8 VSS 0.0046183f
c5 9 VSS 0.0245824f
r1 21 20 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r2 7 20 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r3 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0540 $Y2=0.2340
r4 18 19 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.2340 $X2=0.0930 $Y2=0.2340
r5 16 19 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1515
+ $Y=0.2340 $X2=0.0930 $Y2=0.2340
r6 9 14 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2205
+ $Y=0.2340 $X2=0.2700 $Y2=0.2340
r7 9 16 16.0901 $w=1.3e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.2205
+ $Y=0.2340 $X2=0.1515 $Y2=0.2340
r8 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2700 $Y2=0.2340
r9 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r10 2 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r11 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r12 12 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r13 1 7 1e-05
.ends

.subckt PM_MAJx3_ASAP7_75t_R%Y VSS 32 26 27 41 44 45 47 13 3 15 17 1 19 2 16 14
c1 1 VSS 0.0105672f
c2 2 VSS 0.0109757f
c3 3 VSS 0.00808504f
c4 4 VSS 0.00799129f
c5 13 VSS 0.00454228f
c6 14 VSS 0.00346591f
c7 15 VSS 0.00451775f
c8 16 VSS 0.00345696f
c9 17 VSS 0.00905148f
c10 18 VSS 0.0104069f
c11 19 VSS 0.00499769f
c12 20 VSS 0.00398178f
c13 21 VSS 0.00425418f
c14 22 VSS 0.00243233f
c15 23 VSS 0.00211112f
r1 16 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4840 $Y2=0.2025
r2 47 16 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r3 45 43 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r4 2 43 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.2025 $X2=0.3925 $Y2=0.2025
r5 15 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r6 44 15 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3635 $Y2=0.2025
r7 4 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.2340
r8 2 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.2025
+ $X2=0.3775 $Y2=0.2340
r9 14 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4840 $Y2=0.0675
r10 41 14 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
r11 21 23 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.2340 $X2=0.4590 $Y2=0.2340
r12 18 36 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r13 18 38 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.2340 $X2=0.3775 $Y2=0.2340
r14 3 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0360
r15 23 35 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r16 23 36 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4185 $Y2=0.2340
r17 20 22 5.11582 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r18 34 35 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1780 $X2=0.4590 $Y2=0.2160
r19 33 34 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1485 $X2=0.4590 $Y2=0.1780
r20 32 33 0.23319 $w=1.3e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1485
r21 32 31 9.91056 $w=1.3e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1475 $X2=0.4590 $Y2=0.1050
r22 19 22 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r23 19 31 11.8927 $w=1.3e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.1050
r24 22 30 8.26388 $w=1.41111e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.0360 $X2=0.4185 $Y2=0.0360
r25 29 30 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3865
+ $Y=0.0360 $X2=0.4185 $Y2=0.0360
r26 28 29 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3775
+ $Y=0.0360 $X2=0.3865 $Y2=0.0360
r27 17 28 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3665
+ $Y=0.0360 $X2=0.3775 $Y2=0.0360
r28 1 28 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3775 $Y2=0.0360
r29 27 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r30 1 25 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r31 13 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r32 26 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
.ends

.subckt PM_MAJx3_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00565509f
.ends

.subckt PM_MAJx3_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.00580102f
.ends

.subckt PM_MAJx3_ASAP7_75t_R%B VSS 22 5 6 7 13 11 1 8 9 2 10 14 12
c1 1 VSS 0.0033074f
c2 2 VSS 0.00669407f
c3 5 VSS 0.00782861f
c4 6 VSS 0.0817923f
c5 7 VSS 0.00201208f
c6 8 VSS 0.00228167f
c7 9 VSS 0.00475285f
c8 10 VSS 0.0030127f
c9 11 VSS 0.00174086f
c10 12 VSS 0.00204196f
c11 13 VSS 0.00187732f
c12 14 VSS 0.00261291f
c13 15 VSS 0.0040392f
r1 1 29 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r2 5 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r3 29 30 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1620 $Y2=0.1350
r4 7 29 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1245
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r5 11 28 2.78149 $w=1.76421e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1890 $Y2=0.1540
r6 11 30 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r7 8 12 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1765 $X2=0.1890 $Y2=0.1980
r8 8 28 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1765 $X2=0.1890 $Y2=0.1540
r9 12 27 4.64701 $w=1.46667e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1980 $X2=0.2160 $Y2=0.1980
r10 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r11 25 26 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2675
+ $Y=0.1980 $X2=0.2430 $Y2=0.1980
r12 24 25 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.1980 $X2=0.2675 $Y2=0.1980
r13 22 23 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M1 $thickness=3.6e-08 $X=0.2890
+ $Y=0.1980 $X2=0.3022 $Y2=0.1980
r14 22 9 0.641272 $w=1.3e-08 $l=2.8e-09 $layer=M1 $thickness=3.6e-08 $X=0.2890
+ $Y=0.1980 $X2=0.2862 $Y2=0.1980
r15 9 24 0.641272 $w=1.3e-08 $l=2.7e-09 $layer=M1 $thickness=3.6e-08 $X=0.2862
+ $Y=0.1980 $X2=0.2835 $Y2=0.1980
r16 15 21 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.3240 $Y2=0.1765
r17 15 23 3.42276 $w=1.5069e-08 $l=2.18e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1980 $X2=0.3022 $Y2=0.1980
r18 20 21 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1565 $X2=0.3240 $Y2=0.1765
r19 10 14 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1465 $X2=0.3240 $Y2=0.1350
r20 10 20 2.3319 $w=1.3e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.1465 $X2=0.3240 $Y2=0.1565
r21 14 18 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3105 $Y2=0.1350
r22 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3105 $Y2=0.1350
r23 13 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2855
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r24 6 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r25 2 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1350
+ $X2=0.2970 $Y2=0.1350
.ends

.subckt PM_MAJx3_ASAP7_75t_R%A VSS 7 3 1 4
c1 1 VSS 0.00819199f
c2 3 VSS 0.00848611f
c3 4 VSS 0.0044334f
r1 7 8 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1160 $X2=0.0810 $Y2=0.1212
r2 4 8 3.20636 $w=1.3e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1212
r3 3 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r4 1 4 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
.ends

.subckt PM_MAJx3_ASAP7_75t_R%NET1 VSS 11 18 19 7 1 2 8 9
c1 1 VSS 0.00531367f
c2 2 VSS 0.0100517f
c3 7 VSS 0.00262896f
c4 8 VSS 0.00459803f
c5 9 VSS 0.0228183f
r1 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 2 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r4 18 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r5 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r6 13 14 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.1620
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r7 12 13 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.0540
+ $Y=0.0360 $X2=0.1620 $Y2=0.0360
r8 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r9 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0540 $Y2=0.0360
r10 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r11 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r12 1 7 1e-05
.ends

.subckt PM_MAJx3_ASAP7_75t_R%MAJI VSS 9 10 11 58 59 70 71 13 3 4 16 15 14 12 1
+ 17 18 19 20
c1 1 VSS 0.0125108f
c2 3 VSS 0.00349526f
c3 4 VSS 0.00373031f
c4 9 VSS 0.0807201f
c5 10 VSS 0.080159f
c6 11 VSS 0.0798296f
c7 12 VSS 0.00630253f
c8 13 VSS 0.00637597f
c9 14 VSS 0.00655122f
c10 15 VSS 0.0109734f
c11 16 VSS 0.00209821f
c12 17 VSS 0.00227645f
c13 18 VSS 0.00228981f
c14 19 VSS 0.00228324f
c15 20 VSS 0.000520834f
r1 71 69 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r2 4 69 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2025 $X2=0.1225 $Y2=0.2025
r3 13 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1080 $Y2=0.2025
r4 70 13 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r5 4 65 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1090 $Y2=0.1980
r6 64 65 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.1980 $X2=0.1090 $Y2=0.1980
r7 63 64 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1980 $X2=0.0950 $Y2=0.1980
r8 62 63 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0565
+ $Y=0.1980 $X2=0.0810 $Y2=0.1980
r9 16 19 1.03257 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0385 $Y=0.1980 $X2=0.0270 $Y2=0.1980
r10 16 62 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0385
+ $Y=0.1980 $X2=0.0565 $Y2=0.1980
r11 19 61 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1980 $X2=0.0270 $Y2=0.1765
r12 60 61 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1350 $X2=0.0270 $Y2=0.1765
r13 14 18 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0935 $X2=0.0270 $Y2=0.0720
r14 14 60 9.67737 $w=1.3e-08 $l=4.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0935 $X2=0.0270 $Y2=0.1350
r15 59 57 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r16 3 57 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.0675 $X2=0.1225 $Y2=0.0675
r17 12 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r18 58 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r19 18 55 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0720 $X2=0.0380 $Y2=0.0720
r20 3 51 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1090 $Y2=0.0720
r21 54 55 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0560
+ $Y=0.0720 $X2=0.0380 $Y2=0.0720
r22 53 54 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0720 $X2=0.0560 $Y2=0.0720
r23 51 52 2.44849 $w=1.3e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1090
+ $Y=0.0720 $X2=0.1195 $Y2=0.0720
r24 50 51 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.0720 $X2=0.1090 $Y2=0.0720
r25 50 53 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0950
+ $Y=0.0720 $X2=0.0810 $Y2=0.0720
r26 49 52 9.32759 $w=1.3e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1595
+ $Y=0.0720 $X2=0.1195 $Y2=0.0720
r27 48 49 13.1752 $w=1.3e-08 $l=5.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0720 $X2=0.1595 $Y2=0.0720
r28 47 48 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.0720 $X2=0.2160 $Y2=0.0720
r29 46 47 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.2675
+ $Y=0.0720 $X2=0.2430 $Y2=0.0720
r30 45 46 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2835
+ $Y=0.0720 $X2=0.2675 $Y2=0.0720
r31 44 45 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.2995
+ $Y=0.0720 $X2=0.2835 $Y2=0.0720
r32 43 44 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3240
+ $Y=0.0720 $X2=0.2995 $Y2=0.0720
r33 42 43 5.71315 $w=1.3e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.3485
+ $Y=0.0720 $X2=0.3240 $Y2=0.0720
r34 15 20 0.915974 $w=1.70909e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3660 $Y=0.0720 $X2=0.3770 $Y2=0.0720
r35 15 42 4.08082 $w=1.3e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.3660
+ $Y=0.0720 $X2=0.3485 $Y2=0.0720
r36 20 39 3.36447 $w=1.71023e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3770 $Y=0.0720 $X2=0.3770 $Y2=0.0935
r37 11 35 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r38 10 29 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r39 17 37 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.3770
+ $Y=0.1160 $X2=0.3770 $Y2=0.1350
r40 17 39 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3770
+ $Y=0.1160 $X2=0.3770 $Y2=0.0935
r41 33 35 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4465 $Y=0.1350 $X2=0.4590 $Y2=0.1350
r42 32 33 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4320 $Y=0.1350 $X2=0.4465 $Y2=0.1350
r43 30 32 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4175 $Y=0.1350 $X2=0.4320 $Y2=0.1350
r44 29 30 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.4050 $Y=0.1350 $X2=0.4175 $Y2=0.1350
r45 27 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3925 $Y=0.1350 $X2=0.4050 $Y2=0.1350
r46 26 27 2.65825 $w=1.53e-08 $l=4.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3880 $Y=0.1350 $X2=0.3925 $Y2=0.1350
r47 25 26 6.49795 $w=1.53e-08 $l=1.1e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3770 $Y=0.1350 $X2=0.3880 $Y2=0.1350
r48 25 37 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3770 $Y=0.1350
+ $X2=0.3770 $Y2=0.1350
r49 24 25 5.90723 $w=1.53e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.3670
+ $Y=0.1350 $X2=0.3770 $Y2=0.1350
r50 23 24 2.06753 $w=1.53e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3635 $Y=0.1350 $X2=0.3670 $Y2=0.1350
r51 9 1 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r52 1 22 2.90696 $w=2.1681e-08 $l=1.05e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r53 1 23 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
r54 9 22 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.3510 $Y=0.1350 $X2=0.3405 $Y2=0.1350
r55 9 23 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.3510 $Y=0.1350 $X2=0.3635 $Y2=0.1350
.ends


*
.SUBCKT MAJx3_ASAP7_75t_R VSS VDD A B C Y
*
* VSS VSS
* VDD VDD
* A A
* B B
* C C
* Y Y
*
*

MM0 N_MM0_d N_MM0_g N_MM0_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM3 N_MM3_d N_MM3_g N_MM3_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM9_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM7_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM6_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 N_MM10_d N_MM11_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@3 N_MM10@3_d N_MM11@3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10@2 N_MM10@2_d N_MM11@2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM0_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM3_g N_MM8_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM11_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@3 N_MM11@3_d N_MM11@3_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11@2 N_MM11@2_d N_MM11@2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "MAJx3_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "MAJx3_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_MAJx3_ASAP7_75t_R%NET17 VSS N_MM3_s N_MM4_d N_NET17_1
+ PM_MAJx3_ASAP7_75t_R%NET17
cc_1 N_NET17_1 N_MM3_g 0.0172305f
cc_2 N_NET17_1 N_MM9_g 0.017434f
x_PM_MAJx3_ASAP7_75t_R%NET16 VSS N_MM9_d N_MM8_s N_NET16_1
+ PM_MAJx3_ASAP7_75t_R%NET16
cc_3 N_NET16_1 N_MM3_g 0.0172841f
cc_4 N_NET16_1 N_MM9_g 0.0174499f
x_PM_MAJx3_ASAP7_75t_R%C VSS C N_MM9_g N_MM7_g N_C_5 N_C_1
+ PM_MAJx3_ASAP7_75t_R%C
cc_5 N_MM9_g N_B_13 0.000633092f
cc_6 N_C_5 N_B_11 0.000682114f
cc_7 N_C_1 N_B_1 0.000688856f
cc_8 N_C_5 N_B_8 0.000774008f
cc_9 N_C_5 N_B_9 0.00127049f
cc_10 N_C_1 N_B_11 0.00206432f
cc_11 N_MM7_g N_MM6_g 0.00336639f
cc_12 N_C_5 N_B_13 0.00353333f
cc_13 N_MM9_g N_MM3_g 0.00826898f
x_PM_MAJx3_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_MAJx3_ASAP7_75t_R%noxref_15
cc_14 N_noxref_15_1 N_MM11@2_g 0.00146547f
cc_15 N_noxref_15_1 N_Y_16 0.0371788f
cc_16 N_noxref_15_1 N_noxref_14_1 0.00179172f
x_PM_MAJx3_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_MAJx3_ASAP7_75t_R%noxref_14
cc_17 N_noxref_14_1 N_MM11@2_g 0.00146849f
cc_18 N_noxref_14_1 N_Y_14 0.037444f
x_PM_MAJx3_ASAP7_75t_R%NET3 VSS N_MM7_d N_MM6_d N_MM5_s N_NET3_7 N_NET3_1
+ N_NET3_2 N_NET3_8 N_NET3_9 PM_MAJx3_ASAP7_75t_R%NET3
cc_19 N_NET3_7 N_A_1 0.000719175f
cc_20 N_NET3_1 N_MM0_g 0.00101396f
cc_21 N_NET3_7 N_MM0_g 0.0343426f
cc_22 N_NET3_2 N_MM6_g 0.00217179f
cc_23 N_NET3_8 N_B_2 0.000724851f
cc_24 N_NET3_9 N_B_9 0.00413213f
cc_25 N_NET3_9 N_B_12 0.0059912f
cc_26 N_NET3_8 N_MM6_g 0.0348943f
cc_27 N_NET3_2 N_MM7_g 0.000942381f
cc_28 N_NET3_8 N_MM7_g 0.0351714f
cc_29 N_NET3_9 N_MAJI_4 0.000494161f
cc_30 N_NET3_9 N_MAJI_13 0.000596436f
cc_31 N_NET3_9 N_MAJI_19 0.000620229f
cc_32 N_NET3_1 N_MAJI_16 0.0006221f
cc_33 N_NET3_7 N_MAJI_13 0.000678968f
cc_34 N_NET3_1 N_MAJI_14 0.000694647f
cc_35 N_NET3_1 N_MAJI_4 0.00409434f
cc_36 N_NET3_9 N_MAJI_16 0.00842228f
x_PM_MAJx3_ASAP7_75t_R%Y VSS Y N_MM10_d N_MM10@3_d N_MM10@2_d N_MM11_d
+ N_MM11@3_d N_MM11@2_d N_Y_13 N_Y_3 N_Y_15 N_Y_17 N_Y_1 N_Y_19 N_Y_2 N_Y_16
+ N_Y_14 PM_MAJx3_ASAP7_75t_R%Y
cc_37 N_Y_13 N_MAJI_20 0.000393906f
cc_38 N_Y_13 N_MM11@2_g 0.00169782f
cc_39 N_Y_13 N_MAJI_1 0.000773193f
cc_40 N_Y_3 N_MM11@2_g 0.000852749f
cc_41 N_Y_15 N_MM11@3_g 0.0307581f
cc_42 N_Y_17 N_MAJI_15 0.00123351f
cc_43 N_Y_1 N_MAJI_17 0.00168433f
cc_44 N_Y_19 N_MAJI_1 0.00198398f
cc_45 N_Y_2 N_MM11@3_g 0.00202115f
cc_46 N_Y_1 N_MM11@3_g 0.0026299f
cc_47 N_Y_17 N_MAJI_20 0.0032707f
cc_48 N_Y_16 N_MM11@2_g 0.0148119f
cc_49 N_Y_15 N_MAJI_1 0.0068021f
cc_50 N_Y_14 N_MM11@2_g 0.0523994f
cc_51 N_Y_13 N_MM11_g 0.0369725f
cc_52 N_Y_13 N_MM11@3_g 0.0684065f
x_PM_MAJx3_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_MAJx3_ASAP7_75t_R%noxref_12
cc_53 N_noxref_12_1 N_MM0_g 0.00144276f
cc_54 N_noxref_12_1 N_MAJI_12 0.000743695f
cc_55 N_noxref_12_1 N_NET1_7 0.0363128f
cc_56 N_noxref_12_1 N_NET3_7 0.00047078f
x_PM_MAJx3_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_MAJx3_ASAP7_75t_R%noxref_13
cc_57 N_noxref_13_1 N_MM0_g 0.00144608f
cc_58 N_noxref_13_1 N_MAJI_13 0.000745819f
cc_59 N_noxref_13_1 N_NET1_7 0.000471978f
cc_60 N_noxref_13_1 N_NET3_7 0.0362063f
cc_61 N_noxref_13_1 N_noxref_12_1 0.00176895f
x_PM_MAJx3_ASAP7_75t_R%B VSS B N_MM3_g N_MM6_g N_B_7 N_B_13 N_B_11 N_B_1 N_B_8
+ N_B_9 N_B_2 N_B_10 N_B_14 N_B_12 PM_MAJx3_ASAP7_75t_R%B
cc_62 N_MM3_g N_A_1 0.00087229f
cc_63 N_B_7 N_A_4 0.00173234f
cc_64 N_MM3_g N_MM0_g 0.00418748f
x_PM_MAJx3_ASAP7_75t_R%A VSS A N_MM0_g N_A_1 N_A_4 PM_MAJx3_ASAP7_75t_R%A
x_PM_MAJx3_ASAP7_75t_R%NET1 VSS N_MM0_s N_MM2_d N_MM1_d N_NET1_7 N_NET1_1
+ N_NET1_2 N_NET1_8 N_NET1_9 PM_MAJx3_ASAP7_75t_R%NET1
cc_65 N_NET1_7 N_A_1 0.000764802f
cc_66 N_NET1_1 N_MM0_g 0.0010127f
cc_67 N_NET1_7 N_MM0_g 0.03441f
cc_68 N_NET1_2 N_MM6_g 0.000891958f
cc_69 N_NET1_8 N_MM6_g 0.0354115f
cc_70 N_NET1_2 N_MM7_g 0.000935143f
cc_71 N_NET1_8 N_MM7_g 0.0352709f
cc_72 N_NET1_7 N_MAJI_12 0.00126889f
cc_73 N_NET1_9 N_MAJI_18 0.00063802f
cc_74 N_NET1_1 N_MAJI_14 0.000681207f
cc_75 N_NET1_2 N_MAJI_15 0.000766633f
cc_76 N_NET1_1 N_MAJI_3 0.00412368f
cc_77 N_NET1_9 N_MAJI_15 0.0222575f
x_PM_MAJx3_ASAP7_75t_R%MAJI VSS N_MM11_g N_MM11@3_g N_MM11@2_g N_MM0_d N_MM3_d
+ N_MM5_d N_MM8_d N_MAJI_13 N_MAJI_3 N_MAJI_4 N_MAJI_16 N_MAJI_15 N_MAJI_14
+ N_MAJI_12 N_MAJI_1 N_MAJI_17 N_MAJI_18 N_MAJI_19 N_MAJI_20
+ PM_MAJx3_ASAP7_75t_R%MAJI
cc_78 N_MAJI_13 N_MM0_g 0.015559f
cc_79 N_MAJI_3 N_MM0_g 0.000910145f
cc_80 N_MAJI_4 N_MM0_g 0.000914101f
cc_81 N_MAJI_3 N_A_1 0.00100546f
cc_82 N_MAJI_16 N_A_4 0.00112121f
cc_83 N_MAJI_15 N_A_4 0.00122683f
cc_84 N_MAJI_13 N_A_1 0.00160354f
cc_85 N_MAJI_14 N_A_4 0.00487662f
cc_86 N_MAJI_12 N_MM0_g 0.0539357f
cc_87 N_MAJI_16 N_MM3_g 0.00055638f
cc_88 N_MAJI_4 N_MM3_g 0.00149095f
cc_89 N_MAJI_1 N_MM3_g 0.000602993f
cc_90 N_MAJI_1 N_B_2 0.00040015f
cc_91 N_MAJI_15 N_B_13 0.000457344f
cc_92 N_MAJI_13 N_MM3_g 0.0158856f
cc_93 N_MAJI_16 N_B_7 0.000645397f
cc_94 N_MAJI_17 N_B_10 0.000657315f
cc_95 N_MAJI_1 N_B_14 0.000713649f
cc_96 N_MAJI_3 N_B_1 0.000846912f
cc_97 N_MAJI_3 N_MM3_g 0.00117149f
cc_98 N_MAJI_15 N_B_14 0.00155771f
cc_99 N_MAJI_15 N_B_7 0.00164709f
cc_100 N_MAJI_17 N_B_14 0.00167571f
cc_101 N_MAJI_13 N_B_1 0.00179921f
cc_102 N_MM11_g N_MM6_g 0.00332484f
cc_103 N_MAJI_15 N_B_11 0.00382598f
cc_104 N_MAJI_12 N_MM3_g 0.055342f
cc_105 N_MAJI_3 N_C_5 0.000148788f
cc_106 N_MAJI_12 N_C_5 0.000517854f
cc_107 N_MAJI_15 N_C_5 0.00410043f
*END of MAJx3_ASAP7_75t_R.pxi
.ENDS
** Design:	FAx1_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "FAx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "FAx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_FAx1_ASAP7_75t_R%noxref_21 VSS 1
c1 1 VSS 0.0429241f
.ends

.subckt PM_FAx1_ASAP7_75t_R%noxref_20 VSS 1
c1 1 VSS 0.0429317f
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET027 VSS 12 13 27 28 8 9 2 7 1
c1 1 VSS 0.00678789f
c2 2 VSS 0.00976364f
c3 7 VSS 0.00333418f
c4 8 VSS 0.00460051f
c5 9 VSS 0.0146458f
r1 28 26 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r2 2 26 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.2025 $X2=0.6625 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.2025 $X2=0.6480 $Y2=0.2025
r4 27 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.2025 $X2=0.6335 $Y2=0.2025
r5 2 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.2025
+ $X2=0.6480 $Y2=0.2340
r6 22 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.2340 $X2=0.6480 $Y2=0.2340
r7 21 22 4.6638 $w=1.3e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.6145
+ $Y=0.2340 $X2=0.6345 $Y2=0.2340
r8 20 21 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5930
+ $Y=0.2340 $X2=0.6145 $Y2=0.2340
r9 19 20 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5815
+ $Y=0.2340 $X2=0.5930 $Y2=0.2340
r10 18 19 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.2340 $X2=0.5815 $Y2=0.2340
r11 17 18 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5535
+ $Y=0.2340 $X2=0.5670 $Y2=0.2340
r12 16 17 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5460
+ $Y=0.2340 $X2=0.5535 $Y2=0.2340
r13 9 16 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.5380
+ $Y=0.2340 $X2=0.5460 $Y2=0.2340
r14 1 9 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.2025
+ $X2=0.5380 $Y2=0.2340
r15 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r16 1 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.2025 $X2=0.5545 $Y2=0.2025
r17 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.2025 $X2=0.5400 $Y2=0.2025
r18 12 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.2025 $X2=0.5255 $Y2=0.2025
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET27 VSS 11 26 27 7 9 1 8 2
c1 1 VSS 0.00821341f
c2 2 VSS 0.00777697f
c3 7 VSS 0.00392751f
c4 8 VSS 0.00337154f
c5 9 VSS 0.0229487f
r1 27 25 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 2 25 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.2025 $X2=0.2700 $Y2=0.2025
r4 26 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.2025 $X2=0.2555 $Y2=0.2025
r5 2 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2025
+ $X2=0.2710 $Y2=0.2340
r6 20 21 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2620
+ $Y=0.2340 $X2=0.2710 $Y2=0.2340
r7 19 20 1.28254 $w=1.3e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.2565
+ $Y=0.2340 $X2=0.2620 $Y2=0.2340
r8 18 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.2340 $X2=0.2565 $Y2=0.2340
r9 17 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.2320
+ $Y=0.2340 $X2=0.2430 $Y2=0.2340
r10 16 17 12.8254 $w=1.3e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1770
+ $Y=0.2340 $X2=0.2320 $Y2=0.2340
r11 15 16 16.3233 $w=1.3e-08 $l=7e-08 $layer=M1 $thickness=3.6e-08 $X=0.1070
+ $Y=0.2340 $X2=0.1770 $Y2=0.2340
r12 14 15 7.11229 $w=1.3e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0765
+ $Y=0.2340 $X2=0.1070 $Y2=0.2340
r13 13 14 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.2340 $X2=0.0765 $Y2=0.2340
r14 12 13 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0520
+ $Y=0.2340 $X2=0.0610 $Y2=0.2340
r15 9 12 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.2340 $X2=0.0520 $Y2=0.2340
r16 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2025
+ $X2=0.0520 $Y2=0.2340
r17 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r18 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2025 $X2=0.0685 $Y2=0.2025
r19 1 7 1e-05
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET25 VSS 11 23 24 7 9 1 8 2
c1 1 VSS 0.0082303f
c2 2 VSS 0.00801658f
c3 7 VSS 0.00395749f
c4 8 VSS 0.00338264f
c5 9 VSS 0.0240914f
r1 24 22 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r2 2 22 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2700 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2555 $Y=0.0675 $X2=0.2700 $Y2=0.0675
r4 23 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2530 $Y=0.0675 $X2=0.2555 $Y2=0.0675
r5 2 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r6 17 18 18.0722 $w=1.3e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.1925
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r7 16 17 19.9377 $w=1.3e-08 $l=8.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1070
+ $Y=0.0360 $X2=0.1925 $Y2=0.0360
r8 15 16 6.06293 $w=1.3e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0360 $X2=0.1070 $Y2=0.0360
r9 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0360 $X2=0.0810 $Y2=0.0360
r10 13 14 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0610
+ $Y=0.0360 $X2=0.0675 $Y2=0.0360
r11 12 13 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.0520
+ $Y=0.0360 $X2=0.0610 $Y2=0.0360
r12 9 12 2.2153 $w=1.3e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0425
+ $Y=0.0360 $X2=0.0520 $Y2=0.0360
r13 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0675
+ $X2=0.0520 $Y2=0.0360
r14 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r15 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0675 $X2=0.0685 $Y2=0.0675
r16 1 7 1e-05
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET067 VSS 12 13 28 29 8 2 7 9 1
c1 1 VSS 0.00715334f
c2 2 VSS 0.0103033f
c3 7 VSS 0.00333123f
c4 8 VSS 0.00463593f
c5 9 VSS 0.0139677f
r1 29 27 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5570 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r2 1 27 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5400 $Y=0.0675 $X2=0.5545 $Y2=0.0675
r3 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.5255 $Y=0.0675 $X2=0.5400 $Y2=0.0675
r4 28 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5230 $Y=0.0675 $X2=0.5255 $Y2=0.0675
r5 1 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.5400 $Y=0.0675
+ $X2=0.5380 $Y2=0.0360
r6 21 22 1.74892 $w=1.3e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.5460
+ $Y=0.0360 $X2=0.5535 $Y2=0.0360
r7 21 23 1.86552 $w=1.3e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.5460
+ $Y=0.0360 $X2=0.5380 $Y2=0.0360
r8 20 22 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.0360 $X2=0.5535 $Y2=0.0360
r9 19 20 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.5815
+ $Y=0.0360 $X2=0.5670 $Y2=0.0360
r10 18 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.5930
+ $Y=0.0360 $X2=0.5815 $Y2=0.0360
r11 17 18 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.6055
+ $Y=0.0360 $X2=0.5930 $Y2=0.0360
r12 16 17 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.0360 $X2=0.6055 $Y2=0.0360
r13 9 14 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.0360 $X2=0.6480 $Y2=0.0360
r14 9 16 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.6345
+ $Y=0.0360 $X2=0.6210 $Y2=0.0360
r15 2 14 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.6480 $Y=0.0675
+ $X2=0.6480 $Y2=0.0360
r16 13 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6650 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r17 2 11 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6480 $Y=0.0675 $X2=0.6625 $Y2=0.0675
r18 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6335 $Y=0.0675 $X2=0.6480 $Y2=0.0675
r19 12 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.6310 $Y=0.0675 $X2=0.6335 $Y2=0.0675
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET36 VSS 2 3 1
c1 1 VSS 0.000998966f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1620 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.0675 $X2=0.1620 $Y2=0.0675
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET079 VSS 2 3 1
c1 1 VSS 0.00096155f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3780 $Y2=0.0675
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET080 VSS 2 3 1
c1 1 VSS 0.000977271f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4320 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.0675 $X2=0.4320 $Y2=0.0675
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET37 VSS 2 3 1
c1 1 VSS 0.00103911f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.2025 $X2=0.1620 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1790 $Y=0.2025 $X2=0.1620 $Y2=0.2025
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET081 VSS 2 3 1
c1 1 VSS 0.000956629f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4320 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4490 $Y=0.2025 $X2=0.4320 $Y2=0.2025
.ends

.subckt PM_FAx1_ASAP7_75t_R%NET082 VSS 2 3 1
c1 1 VSS 0.000947645f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.2025 $X2=0.3780 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.2025 $X2=0.3780 $Y2=0.2025
.ends

.subckt PM_FAx1_ASAP7_75t_R%noxref_18 VSS 1
c1 1 VSS 0.00603683f
.ends

.subckt PM_FAx1_ASAP7_75t_R%noxref_19 VSS 1
c1 1 VSS 0.00606537f
.ends

.subckt PM_FAx1_ASAP7_75t_R%SN VSS 39 19 20 50 51 11 9 10 8 12 7 1 2 15 16
c1 1 VSS 0.00380077f
c2 2 VSS 0.00348579f
c3 7 VSS 0.00242227f
c4 8 VSS 0.00242675f
c5 9 VSS 0.00593461f
c6 10 VSS 0.0123256f
c7 11 VSS 0.012642f
c8 12 VSS 0.000461433f
c9 13 VSS 0.00361295f
c10 14 VSS 0.00375138f
c11 15 VSS 0.00254304f
c12 16 VSS 0.00204051f
r1 51 49 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r2 2 49 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.2025 $X2=0.5005 $Y2=0.2025
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.2025 $X2=0.4860 $Y2=0.2025
r4 50 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.2025 $X2=0.4715 $Y2=0.2025
r5 2 47 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.2025
+ $X2=0.4860 $Y2=0.1935
r6 12 45 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2025 $X2=0.4860 $Y2=0.2160
r7 12 47 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2025 $X2=0.4860 $Y2=0.1935
r8 16 44 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4860 $Y=0.2340 $X2=0.4725 $Y2=0.2340
r9 16 45 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.2340 $X2=0.4860 $Y2=0.2160
r10 43 44 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4725 $Y2=0.2340
r11 42 43 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4590 $Y2=0.2340
r12 41 42 7.81186 $w=1.3e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3985
+ $Y=0.2340 $X2=0.4320 $Y2=0.2340
r13 11 14 5.22999 $w=1.45254e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3625 $Y=0.2340 $X2=0.3330 $Y2=0.2340
r14 11 41 8.39483 $w=1.3e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.3625
+ $Y=0.2340 $X2=0.3985 $Y2=0.2340
r15 14 40 1.55725 $w=1.94145e-08 $l=1.38e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3330 $Y=0.2340 $X2=0.3330 $Y2=0.2202
r16 39 40 1.22425 $w=1.3e-08 $l=5.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.2150 $X2=0.3330 $Y2=0.2202
r17 39 38 0.991057 $w=1.3e-08 $l=4.3e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.2150 $X2=0.3330 $Y2=0.2107
r18 37 38 1.92382 $w=1.3e-08 $l=8.2e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.2025 $X2=0.3330 $Y2=0.2107
r19 36 37 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1935 $X2=0.3330 $Y2=0.2025
r20 35 36 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1845 $X2=0.3330 $Y2=0.1935
r21 34 35 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1735 $X2=0.3330 $Y2=0.1845
r22 33 34 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1440 $X2=0.3330 $Y2=0.1735
r23 32 33 6.8791 $w=1.3e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1145 $X2=0.3330 $Y2=0.1440
r24 31 32 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.1055 $X2=0.3330 $Y2=0.1145
r25 30 31 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.0965 $X2=0.3330 $Y2=0.1055
r26 29 30 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.0810 $X2=0.3330 $Y2=0.0965
r27 28 29 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.0700 $X2=0.3330 $Y2=0.0810
r28 9 13 3.13128 $w=1.73024e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3330 $Y=0.0565 $X2=0.3330 $Y2=0.0360
r29 9 28 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3330
+ $Y=0.0565 $X2=0.3330 $Y2=0.0700
r30 13 27 5.22999 $w=1.45254e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3330 $Y=0.0360 $X2=0.3625 $Y2=0.0360
r31 26 27 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.3895
+ $Y=0.0360 $X2=0.3625 $Y2=0.0360
r32 25 26 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.0360 $X2=0.3895 $Y2=0.0360
r33 24 25 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4050 $Y2=0.0360
r34 23 24 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0360 $X2=0.4320 $Y2=0.0360
r35 10 22 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4725 $Y=0.0360 $X2=0.4860 $Y2=0.0360
r36 10 23 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4725
+ $Y=0.0360 $X2=0.4590 $Y2=0.0360
r37 15 22 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4860
+ $Y=0.0540 $X2=0.4860 $Y2=0.0360
r38 1 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4860 $Y=0.0675
+ $X2=0.4860 $Y2=0.0540
r39 20 18 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.5030 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r40 1 18 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4860 $Y=0.0675 $X2=0.5005 $Y2=0.0675
r41 7 1 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4715 $Y=0.0675 $X2=0.4860 $Y2=0.0675
r42 19 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4690 $Y=0.0675 $X2=0.4715 $Y2=0.0675
.ends

.subckt PM_FAx1_ASAP7_75t_R%CON VSS 30 9 56 57 67 68 12 10 11 13 3 4 16 17 15
+ 21 14 18 1 20 19
c1 1 VSS 9.22244e-20
c2 3 VSS 0.00359839f
c3 4 VSS 0.00366007f
c4 9 VSS 0.00449162f
c5 10 VSS 0.00508015f
c6 11 VSS 0.00515584f
c7 12 VSS 0.00160811f
c8 13 VSS 0.00133305f
c9 14 VSS 0.000838034f
c10 15 VSS 8.99443e-20
c11 16 VSS 0.000688622f
c12 17 VSS 0.000555696f
c13 18 VSS 6.23308e-20
c14 19 VSS 0.000478091f
c15 20 VSS 0.000231202f
c16 21 VSS 0.0121794f
r1 68 66 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r2 4 66 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.2025 $X2=0.2305 $Y2=0.2025
r3 11 4 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.2025 $X2=0.2160 $Y2=0.2025
r4 67 11 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.2025 $X2=0.2015 $Y2=0.2025
r5 4 62 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.2025
+ $X2=0.2160 $Y2=0.1980
r6 61 62 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.1980 $X2=0.2160 $Y2=0.1980
r7 60 61 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1980 $X2=0.2025 $Y2=0.1980
r8 59 60 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1735
+ $Y=0.1980 $X2=0.1890 $Y2=0.1980
r9 14 17 3.37407 $w=1.43235e-08 $l=2.19659e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1545 $Y=0.1980 $X2=0.1330 $Y2=0.1935
r10 14 59 4.43061 $w=1.3e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1545
+ $Y=0.1980 $X2=0.1735 $Y2=0.1980
r11 17 53 1.50855 $w=1.55e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1935 $X2=0.1330 $Y2=0.1845
r12 57 55 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2330 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r13 3 55 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2160 $Y=0.0675 $X2=0.2305 $Y2=0.0675
r14 10 3 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2015 $Y=0.0675 $X2=0.2160 $Y2=0.0675
r15 56 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1990 $Y=0.0675 $X2=0.2015 $Y2=0.0675
r16 52 53 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1735 $X2=0.1330 $Y2=0.1845
r17 51 52 2.09871 $w=1.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1645 $X2=0.1330 $Y2=0.1735
r18 50 51 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1530 $X2=0.1330 $Y2=0.1645
r19 49 50 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1325 $X2=0.1330 $Y2=0.1530
r20 48 49 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.1145 $X2=0.1330 $Y2=0.1325
r21 12 16 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.0990 $X2=0.1330 $Y2=0.0810
r22 12 48 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1330
+ $Y=0.0990 $X2=0.1330 $Y2=0.1145
r23 3 42 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2160 $Y=0.0675
+ $X2=0.2160 $Y2=0.0810
r24 16 36 39.0693 $w=1.8e-08 $l=9e-09 $layer=V1 $X=0.1330 $Y=0.0810 $X2=0.1420
+ $Y2=0.0810
r25 41 42 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.2025
+ $Y=0.0810 $X2=0.2160 $Y2=0.0810
r26 40 41 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.0810 $X2=0.2025 $Y2=0.0810
r27 39 40 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.1735
+ $Y=0.0810 $X2=0.1890 $Y2=0.0810
r28 38 39 3.38125 $w=1.3e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1590
+ $Y=0.0810 $X2=0.1735 $Y2=0.0810
r29 13 38 2.91487 $w=1.3e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1465
+ $Y=0.0810 $X2=0.1590 $Y2=0.0810
r30 13 36 39.0693 $w=1.8e-08 $l=9e-09 $layer=V1 $X=0.1465 $Y=0.0810 $X2=0.1420
+ $Y2=0.0810
r31 13 16 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1465 $Y=0.0810 $X2=0.1330 $Y2=0.0810
r32 36 37 3.96423 $w=1.3e-08 $l=1.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.1420
+ $Y=0.0810 $X2=0.1590 $Y2=0.0810
r33 34 37 9.0944 $w=1.3e-08 $l=3.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.1980
+ $Y=0.0810 $X2=0.1590 $Y2=0.0810
r34 31 32 28.8572 $w=1.3e-08 $l=1.238e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.4052 $Y=0.0810 $X2=0.5290 $Y2=0.0810
r35 30 31 26.8751 $w=1.3e-08 $l=1.152e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2900 $Y=0.0810 $X2=0.4052 $Y2=0.0810
r36 30 21 7.17059 $w=1.3e-08 $l=3.08e-08 $layer=M2 $thickness=3.6e-08 $X=0.2900
+ $Y=0.0810 $X2=0.2592 $Y2=0.0810
r37 21 34 14.2829 $w=1.3e-08 $l=6.12e-08 $layer=M2 $thickness=3.6e-08 $X=0.2592
+ $Y=0.0810 $X2=0.1980 $Y2=0.0810
r38 20 28 1.50137 $w=1.6913e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5355 $Y=0.0810 $X2=0.5240 $Y2=0.0810
r39 20 32 70.3248 $w=1.8e-08 $l=5e-09 $layer=V1 $X=0.5355 $Y=0.0810 $X2=0.5290
+ $Y2=0.0810
r40 28 32 27.048 $w=1.8e-08 $l=1.3e-08 $layer=V1 $X=0.5240 $Y=0.0810 $X2=0.5290
+ $Y2=0.0810
r41 19 27 2.9921 $w=1.50645e-08 $l=1.47139e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5240 $Y=0.0990 $X2=0.5095 $Y2=0.0965
r42 19 28 1.8368 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5240
+ $Y=0.0990 $X2=0.5240 $Y2=0.0810
r43 18 27 2.87127 $w=1.1e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5095
+ $Y=0.1055 $X2=0.5095 $Y2=0.0965
r44 15 25 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5130
+ $Y=0.1170 $X2=0.5130 $Y2=0.1350
r45 15 18 2.89628 $w=1.25652e-08 $l=1.20208e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1170 $X2=0.5095 $Y2=0.1055
r46 15 19 3.01711 $w=1.55e-08 $l=2.1095e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.5130 $Y=0.1170 $X2=0.5240 $Y2=0.0990
r47 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5130
+ $Y=0.1350 $X2=0.5130 $Y2=0.1350
r48 1 25 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5130 $Y=0.1350
+ $X2=0.5130 $Y2=0.1350
.ends

.subckt PM_FAx1_ASAP7_75t_R%CI VSS 23 7 8 9 10 14 15 3 2 16 11 13 1 12
c1 1 VSS 0.00462615f
c2 2 VSS 0.00469392f
c3 3 VSS 0.0080673f
c4 7 VSS 0.00675475f
c5 8 VSS 0.00807732f
c6 9 VSS 0.0822886f
c7 10 VSS 0.00474834f
c8 11 VSS 0.00227199f
c9 12 VSS 0.00458125f
c10 13 VSS 0.00230904f
c11 14 VSS 0.00507295f
c12 15 VSS 0.00268605f
c13 16 VSS 0.00344484f
r1 3 33 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.5670 $Y=0.1350
+ $X2=0.5670 $Y2=0.1350
r2 9 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.5670
+ $Y=0.1350 $X2=0.5670 $Y2=0.1350
r3 2 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4590 $Y=0.1350
+ $X2=0.4590 $Y2=0.1325
r4 8 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4590
+ $Y=0.1350 $X2=0.4590 $Y2=0.1350
r5 15 28 58.604 $w=1.8e-08 $l=6e-09 $layer=V1 $X=0.5790 $Y=0.1170 $X2=0.5730
+ $Y2=0.1170
r6 14 28 29.302 $w=1.8e-08 $l=1.2e-08 $layer=V1 $X=0.5670 $Y=0.1170 $X2=0.5730
+ $Y2=0.1170
r7 14 33 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1170 $X2=0.5670 $Y2=0.1350
r8 14 15 1.61797 $w=1.675e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.5670
+ $Y=0.1170 $X2=0.5790 $Y2=0.1170
r9 10 25 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.4590 $Y=0.1145 $X2=0.4590
+ $Y2=0.1170
r10 10 31 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1145 $X2=0.4590 $Y2=0.1325
r11 27 28 4.5472 $w=1.3e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.5535
+ $Y=0.1170 $X2=0.5730 $Y2=0.1170
r12 26 27 11.1931 $w=1.3e-08 $l=4.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.5055
+ $Y=0.1170 $X2=0.5535 $Y2=0.1170
r13 25 26 10.8433 $w=1.3e-08 $l=4.65e-08 $layer=M2 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1170 $X2=0.5055 $Y2=0.1170
r14 24 25 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1170 $X2=0.4590 $Y2=0.1170
r15 23 24 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1170 $X2=0.3510 $Y2=0.1170
r16 23 16 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1170 $X2=0.2315 $Y2=0.1170
r17 11 12 1.85116 $w=1.64615e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2300 $Y=0.1170 $X2=0.2430 $Y2=0.1170
r18 12 21 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2430
+ $Y=0.1170 $X2=0.2430 $Y2=0.1350
r19 12 13 2.20094 $w=1.61034e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2430 $Y=0.1170 $X2=0.2575 $Y2=0.1170
r20 23 12 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2430 $Y=0.1170
+ $X2=0.2430 $Y2=0.1170
r21 7 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.2430
+ $Y=0.1350 $X2=0.2430 $Y2=0.1350
r22 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2430 $Y=0.1350
+ $X2=0.2430 $Y2=0.1350
.ends

.subckt PM_FAx1_ASAP7_75t_R%B VSS 29 7 8 9 10 14 13 11 15 1 12 2 3
c1 1 VSS 0.00487113f
c2 2 VSS 0.0141572f
c3 3 VSS 0.00887892f
c4 7 VSS 0.00855689f
c5 8 VSS 0.0823298f
c6 9 VSS 0.0854721f
c7 10 VSS 0.0826679f
c8 11 VSS 0.00499223f
c9 12 VSS 0.00683756f
c10 13 VSS 0.0045801f
c11 14 VSS 0.00234643f
c12 15 VSS 0.00487603f
r1 9 46 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r2 8 38 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r3 1 35 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.1890 $Y=0.1350
+ $X2=0.1890 $Y2=0.1350
r4 7 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.1890
+ $Y=0.1350 $X2=0.1890 $Y2=0.1350
r5 44 46 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3385 $Y=0.1350 $X2=0.3510 $Y2=0.1350
r6 43 44 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3240 $Y=0.1350 $X2=0.3385 $Y2=0.1350
r7 41 43 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.3095 $Y=0.1350 $X2=0.3240 $Y2=0.1350
r8 39 41 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.3065 $Y=0.1350 $X2=0.3095 $Y2=0.1350
r9 38 39 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2970
+ $Y=0.1350 $X2=0.3065 $Y2=0.1350
r10 2 38 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.2875
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r11 14 34 1.18787 $w=1.49231e-08 $l=1.45344e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1465 $X2=0.1760 $Y2=0.1530
r12 14 35 2.35382 $w=1.4087e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1890 $Y=0.1465 $X2=0.1890 $Y2=0.1350
r13 14 37 0.9184 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1890
+ $Y=0.1465 $X2=0.1890 $Y2=0.1555
r14 34 37 1.59605 $w=1.60952e-08 $l=1.32382e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1760 $Y=0.1530 $X2=0.1890 $Y2=0.1555
r15 13 34 1.51573 $w=1.3e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1695
+ $Y=0.1530 $X2=0.1760 $Y2=0.1530
r16 11 32 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2970
+ $Y=0.1375 $X2=0.2970 $Y2=0.1555
r17 11 38 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.2970 $Y=0.1375
+ $X2=0.2970 $Y2=0.1350
r18 29 30 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.1810
+ $Y=0.1530 $X2=0.2095 $Y2=0.1530
r19 29 34 43.953 $w=1.8e-08 $l=8e-09 $layer=V1 $X=0.1810 $Y=0.1530 $X2=0.1760
+ $Y2=0.1530
r20 29 37 35.1624 $w=1.8e-08 $l=1e-08 $layer=V1 $X=0.1810 $Y=0.1530 $X2=0.1890
+ $Y2=0.1555
r21 26 27 34.8619 $w=1.3e-08 $l=1.495e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2970 $Y=0.1530 $X2=0.4465 $Y2=0.1530
r22 26 32 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.2970 $Y=0.1530
+ $X2=0.2970 $Y2=0.1555
r23 25 26 8.97781 $w=1.3e-08 $l=3.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1530 $X2=0.2970 $Y2=0.1530
r24 25 30 11.4263 $w=1.3e-08 $l=4.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.2585
+ $Y=0.1530 $X2=0.2095 $Y2=0.1530
r25 24 27 37.427 $w=1.3e-08 $l=1.605e-07 $layer=M2 $thickness=3.6e-08 $X=0.6070
+ $Y=0.1530 $X2=0.4465 $Y2=0.1530
r26 15 22 6.64591 $w=1.3e-08 $l=2.85e-08 $layer=M2 $thickness=3.6e-08 $X=0.6465
+ $Y=0.1530 $X2=0.6750 $Y2=0.1530
r27 15 24 9.211 $w=1.3e-08 $l=3.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.6465
+ $Y=0.1530 $X2=0.6070 $Y2=0.1530
r28 20 22 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6750 $Y=0.1440
+ $X2=0.6750 $Y2=0.1530
r29 12 20 4.78039 $w=1.3e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.6750
+ $Y=0.1235 $X2=0.6750 $Y2=0.1440
r30 10 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.6750
+ $Y=0.1350 $X2=0.6750 $Y2=0.1350
r31 3 20 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6750 $Y=0.1350
+ $X2=0.6750 $Y2=0.1440
.ends

.subckt PM_FAx1_ASAP7_75t_R%A VSS 37 7 8 9 10 17 15 1 16 2 13 12 3 11 14
c1 1 VSS 0.0104824f
c2 2 VSS 0.000812658f
c3 3 VSS 0.00377668f
c4 7 VSS 0.0799284f
c5 8 VSS 0.0828636f
c6 9 VSS 0.00822695f
c7 10 VSS 0.0801077f
c8 11 VSS 0.00351415f
c9 12 VSS 0.000484322f
c10 13 VSS 0.000950982f
c11 14 VSS 0.00335224f
c12 15 VSS 0.000691809f
c13 16 VSS 0.00147063f
c14 17 VSS 0.0371917f
r1 3 49 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.6210 $Y=0.1350
+ $X2=0.6210 $Y2=0.1350
r2 10 3 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1350
r3 2 46 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
r4 9 2 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r5 49 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1350 $X2=0.6210 $Y2=0.1465
r6 48 50 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1580 $X2=0.6210 $Y2=0.1465
r7 13 16 2.02318 $w=2.05484e-08 $l=1.68077e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.6210 $Y=0.1735 $X2=0.6145 $Y2=0.1890
r8 13 48 3.61444 $w=1.3e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.6210
+ $Y=0.1735 $X2=0.6210 $Y2=0.1580
r9 46 47 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1465
r10 12 15 3.72721 $w=1.44857e-08 $l=1.86682e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1645 $X2=0.3985 $Y2=0.1820
r11 12 47 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1645 $X2=0.4050 $Y2=0.1465
r12 16 42 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.6145 $Y=0.1890
+ $X2=0.6130 $Y2=0.1890
r13 15 44 0.507446 $w=2.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.3985
+ $Y=0.1820 $X2=0.3985 $Y2=0.1910
r14 41 42 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.5050
+ $Y=0.1890 $X2=0.6130 $Y2=0.1890
r15 40 41 25.1845 $w=1.3e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.3970
+ $Y=0.1890 $X2=0.5050 $Y2=0.1890
r16 40 44 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.3970 $Y=0.1890
+ $X2=0.3985 $Y2=0.1910
r17 39 40 27.8662 $w=1.3e-08 $l=1.195e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.2775 $Y=0.1890 $X2=0.3970 $Y2=0.1890
r18 38 39 28.7406 $w=1.3e-08 $l=1.233e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.1542 $Y=0.1890 $X2=0.2775 $Y2=0.1890
r19 37 38 3.08976 $w=1.3e-08 $l=1.32e-08 $layer=M2 $thickness=3.6e-08 $X=0.1410
+ $Y=0.1890 $X2=0.1542 $Y2=0.1890
r20 37 36 1.57403 $w=1.3e-08 $l=6.8e-09 $layer=M2 $thickness=3.6e-08 $X=0.1410
+ $Y=0.1890 $X2=0.1342 $Y2=0.1890
r21 35 36 6.8208 $w=1.3e-08 $l=2.92e-08 $layer=M2 $thickness=3.6e-08 $X=0.1050
+ $Y=0.1890 $X2=0.1342 $Y2=0.1890
r22 34 35 7.46207 $w=1.3e-08 $l=3.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.0730
+ $Y=0.1890 $X2=0.1050 $Y2=0.1890
r23 17 34 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M2 $thickness=3.6e-08 $X=0.0615
+ $Y=0.1890 $X2=0.0730 $Y2=0.1890
r24 14 32 4.70486 $w=1.73333e-08 $l=2.77714e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0745 $Y=0.1890 $X2=0.0810 $Y2=0.1620
r25 14 34 19.5347 $w=1.8e-08 $l=1.8e-08 $layer=V1 $X=0.0745 $Y=0.1890
+ $X2=0.0730 $Y2=0.1890
r26 8 29 2.92627 $w=1.245e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r27 31 32 6.29612 $w=1.3e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0810 $Y2=0.1620
r28 11 31 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1235 $X2=0.0810 $Y2=0.1350
r29 27 29 4.08841 $w=2.066e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1225 $Y=0.1350 $X2=0.1350 $Y2=0.1350
r30 26 27 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1080 $Y=0.1350 $X2=0.1225 $Y2=0.1350
r31 25 26 8.56549 $w=1.53e-08 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.0935 $Y=0.1350 $X2=0.1080 $Y2=0.1350
r32 23 25 1.60739 $w=1.64167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0905 $Y=0.1350 $X2=0.0935 $Y2=0.1350
r33 22 23 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1350 $X2=0.0905 $Y2=0.1350
r34 22 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1350
+ $X2=0.0810 $Y2=0.1350
r35 1 22 2.48102 $w=2.2e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0810 $Y2=0.1350
r36 1 24 0.425942 $w=1.865e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.0715
+ $Y=0.1350 $X2=0.0705 $Y2=0.1350
r37 7 22 2.66511 $w=1.29895e-07 $l=0 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0810 $Y2=0.1350
r38 7 24 0.610027 $w=2.16919e-07 $l=1.05e-08 $layer=Gate_1
+ $thickness=5.5619e-08 $X=0.0810 $Y=0.1350 $X2=0.0705 $Y2=0.1350
r39 7 25 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0935 $Y2=0.1350
.ends


*
.SUBCKT FAx1_ASAP7_75t_R VSS VDD A B CI CON SN
*
* VSS VSS
* VDD VDD
* A A
* B B
* CI CI
* CON CON
* SN SN
*
*

MM9 VSS N_MM9_g N_MM9_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM10 VSS N_MM6_g N_MM10_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM8 N_MM8_d N_MM5_g N_MM8_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM7 N_MM7_d N_MM1_g N_MM7_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 VSS N_MM2_g N_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM23 N_MM23_d N_MM20_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM24 N_MM24_d N_MM21_g N_MM24_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM25 N_MM25_d N_MM22_g N_MM25_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM16 N_MM16_d N_MM15_g N_MM16_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM19 VSS N_MM14_g N_MM19_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM17 VSS N_MM17_g N_MM17_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM18 VSS N_MM18_g N_MM18_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g N_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g N_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM20 N_MM20_d N_MM20_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM21 N_MM21_d N_MM21_g N_MM21_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM22 N_MM22_d N_MM22_g N_MM22_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM15 N_MM15_d N_MM15_g N_MM15_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM14 N_MM14_d N_MM14_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM12 N_MM12_d N_MM17_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM13 N_MM13_d N_MM18_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "FAx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "FAx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_FAx1_ASAP7_75t_R%noxref_21 VSS N_noxref_21_1 PM_FAx1_ASAP7_75t_R%noxref_21
cc_1 N_noxref_21_1 N_MM18_g 0.00163289f
cc_2 N_noxref_21_1 N_noxref_20_1 0.00179383f
x_PM_FAx1_ASAP7_75t_R%noxref_20 VSS N_noxref_20_1 PM_FAx1_ASAP7_75t_R%noxref_20
cc_3 N_noxref_20_1 N_MM18_g 0.00163793f
x_PM_FAx1_ASAP7_75t_R%NET027 VSS N_MM15_s N_MM14_d N_MM12_d N_MM13_d N_NET027_8
+ N_NET027_9 N_NET027_2 N_NET027_7 N_NET027_1 PM_FAx1_ASAP7_75t_R%NET027
cc_4 N_NET027_8 N_A_16 0.000462263f
cc_5 N_NET027_8 N_A_3 0.000941512f
cc_6 N_NET027_8 N_A_13 0.000361615f
cc_7 N_NET027_9 N_A_17 0.000830567f
cc_8 N_NET027_2 N_MM17_g 0.0011857f
cc_9 N_NET027_9 N_A_16 0.00362194f
cc_10 N_NET027_8 N_MM17_g 0.0332339f
cc_11 N_NET027_8 N_B_12 0.000376903f
cc_12 N_NET027_8 N_B_3 0.00060497f
cc_13 N_NET027_9 N_B_15 0.000621988f
cc_14 N_NET027_2 N_MM18_g 0.000993449f
cc_15 N_NET027_8 N_MM18_g 0.0333381f
cc_16 N_NET027_7 N_CI_3 0.00103976f
cc_17 N_NET027_1 N_MM14_g 0.000923893f
cc_18 N_NET027_7 N_MM14_g 0.03354f
cc_19 N_NET027_7 N_CON_1 0.00063918f
cc_20 N_NET027_1 N_MM15_g 0.00089605f
cc_21 N_NET027_7 N_MM15_g 0.0335453f
cc_22 N_NET027_7 N_SN_8 0.000557831f
cc_23 N_NET027_9 N_SN_16 0.00101764f
cc_24 N_NET027_1 N_SN_2 0.00442479f
x_PM_FAx1_ASAP7_75t_R%NET27 VSS N_MM0_d N_MM1_s N_MM2_d N_NET27_7 N_NET27_9
+ N_NET27_1 N_NET27_8 N_NET27_2 PM_FAx1_ASAP7_75t_R%NET27
cc_25 N_NET27_7 N_A_1 0.00115805f
cc_26 N_NET27_7 N_A_14 0.000359861f
cc_27 N_NET27_7 N_A_11 0.000392468f
cc_28 N_NET27_9 N_A_14 0.00152646f
cc_29 N_NET27_1 N_MM9_g 0.00161603f
cc_30 N_NET27_9 N_A_17 0.00428946f
cc_31 N_NET27_7 N_MM9_g 0.0341085f
cc_32 N_NET27_8 N_B_15 8.95036e-20
cc_33 N_NET27_8 N_B_2 0.000940744f
cc_34 N_NET27_8 N_B_13 0.000323771f
cc_35 N_NET27_8 N_B_11 0.000355889f
cc_36 N_NET27_2 N_MM2_g 0.00105543f
cc_37 N_NET27_8 N_MM2_g 0.033956f
cc_38 N_NET27_8 N_CI_1 0.000609328f
cc_39 N_NET27_2 N_MM1_g 0.000904302f
cc_40 N_NET27_8 N_MM1_g 0.0340971f
cc_41 N_NET27_9 N_CON_4 0.000816739f
cc_42 N_NET27_9 N_CON_11 0.000561619f
cc_43 N_NET27_8 N_CON_11 0.00058782f
cc_44 N_NET27_9 N_CON_17 0.00082134f
cc_45 N_NET27_2 N_CON_4 0.0030935f
cc_46 N_NET27_9 N_CON_14 0.0088933f
x_PM_FAx1_ASAP7_75t_R%NET25 VSS N_MM9_s N_MM7_d N_MM11_s N_NET25_7 N_NET25_9
+ N_NET25_1 N_NET25_8 N_NET25_2 PM_FAx1_ASAP7_75t_R%NET25
cc_47 N_NET25_7 N_A_17 0.000132631f
cc_48 N_NET25_7 N_A_1 0.00124611f
cc_49 N_NET25_7 N_A_11 0.00044632f
cc_50 N_NET25_9 N_MM6_g 0.00047819f
cc_51 N_NET25_1 N_MM9_g 0.00123352f
cc_52 N_NET25_7 N_MM9_g 0.0340484f
cc_53 N_NET25_8 N_B_14 0.000145695f
cc_54 N_NET25_8 N_B_2 0.000929788f
cc_55 N_NET25_2 N_MM2_g 0.000879282f
cc_56 N_NET25_8 N_MM2_g 0.0339961f
cc_57 N_NET25_8 N_CI_1 0.000716202f
cc_58 N_NET25_2 N_MM1_g 0.000907424f
cc_59 N_NET25_8 N_MM1_g 0.0340884f
cc_60 N_NET25_9 N_CON_3 0.000383174f
cc_61 N_NET25_8 N_CON_10 0.00116674f
cc_62 N_NET25_9 N_CON_16 0.000719495f
cc_63 N_NET25_9 N_CON_21 0.00111465f
cc_64 N_NET25_2 N_CON_3 0.00353584f
cc_65 N_NET25_9 N_CON_13 0.0109273f
x_PM_FAx1_ASAP7_75t_R%NET067 VSS N_MM17_s N_MM18_s N_MM16_d N_MM19_s N_NET067_8
+ N_NET067_2 N_NET067_7 N_NET067_9 N_NET067_1 PM_FAx1_ASAP7_75t_R%NET067
cc_66 N_NET067_8 N_A_13 0.000555978f
cc_67 N_NET067_8 N_A_3 0.000872171f
cc_68 N_NET067_2 N_MM17_g 0.000916733f
cc_69 N_NET067_8 N_MM17_g 0.033206f
cc_70 N_NET067_8 N_B_3 0.000933609f
cc_71 N_NET067_8 N_B_12 0.000661228f
cc_72 N_NET067_2 N_MM18_g 0.000957967f
cc_73 N_NET067_8 N_MM18_g 0.0333647f
cc_74 N_NET067_7 N_CI_3 0.000807629f
cc_75 N_NET067_7 N_CI_14 0.000262354f
cc_76 N_NET067_7 N_CI_15 0.000289238f
cc_77 N_NET067_9 N_CI_15 0.000519807f
cc_78 N_NET067_1 N_MM14_g 0.000924259f
cc_79 N_NET067_7 N_MM14_g 0.0334669f
cc_80 N_NET067_7 N_CON_20 0.000197971f
cc_81 N_NET067_7 N_CON_21 0.000271301f
cc_82 N_NET067_7 N_CON_19 0.000285928f
cc_83 N_NET067_9 N_CON_19 0.000521132f
cc_84 N_NET067_7 N_CON_1 0.000687097f
cc_85 N_NET067_1 N_MM15_g 0.00130249f
cc_86 N_NET067_9 N_CON_20 0.00186215f
cc_87 N_NET067_7 N_MM15_g 0.0335144f
cc_88 N_NET067_9 N_SN_15 0.0010761f
cc_89 N_NET067_1 N_SN_1 0.00435302f
x_PM_FAx1_ASAP7_75t_R%NET36 VSS N_MM10_s N_MM8_d N_NET36_1
+ PM_FAx1_ASAP7_75t_R%NET36
cc_90 N_NET36_1 N_MM6_g 0.0173022f
cc_91 N_NET36_1 N_MM5_g 0.0173474f
x_PM_FAx1_ASAP7_75t_R%NET079 VSS N_MM23_d N_MM24_s N_NET079_1
+ PM_FAx1_ASAP7_75t_R%NET079
cc_92 N_NET079_1 N_MM21_g 0.0173313f
cc_93 N_NET079_1 N_MM20_g 0.0172747f
x_PM_FAx1_ASAP7_75t_R%NET080 VSS N_MM24_d N_MM25_s N_NET080_1
+ PM_FAx1_ASAP7_75t_R%NET080
cc_94 N_NET080_1 N_MM21_g 0.0174102f
cc_95 N_NET080_1 N_MM22_g 0.0171741f
x_PM_FAx1_ASAP7_75t_R%NET37 VSS N_MM6_d N_MM5_s N_NET37_1
+ PM_FAx1_ASAP7_75t_R%NET37
cc_96 N_NET37_1 N_MM6_g 0.0173862f
cc_97 N_NET37_1 N_MM5_g 0.0174368f
x_PM_FAx1_ASAP7_75t_R%NET081 VSS N_MM21_d N_MM22_s N_NET081_1
+ PM_FAx1_ASAP7_75t_R%NET081
cc_98 N_NET081_1 N_MM21_g 0.0174509f
cc_99 N_NET081_1 N_MM22_g 0.0171948f
x_PM_FAx1_ASAP7_75t_R%NET082 VSS N_MM20_d N_MM21_s N_NET082_1
+ PM_FAx1_ASAP7_75t_R%NET082
cc_100 N_NET082_1 N_MM21_g 0.0173746f
cc_101 N_NET082_1 N_MM20_g 0.0172846f
x_PM_FAx1_ASAP7_75t_R%noxref_18 VSS N_noxref_18_1 PM_FAx1_ASAP7_75t_R%noxref_18
cc_102 N_noxref_18_1 N_MM9_g 0.00167063f
cc_103 N_noxref_18_1 N_NET25_7 0.0363075f
cc_104 N_noxref_18_1 N_NET27_7 0.00054419f
x_PM_FAx1_ASAP7_75t_R%noxref_19 VSS N_noxref_19_1 PM_FAx1_ASAP7_75t_R%noxref_19
cc_105 N_noxref_19_1 N_MM9_g 0.00174742f
cc_106 N_noxref_19_1 N_NET25_7 0.000564902f
cc_107 N_noxref_19_1 N_NET27_7 0.0362407f
cc_108 N_noxref_19_1 N_noxref_18_1 0.00179247f
x_PM_FAx1_ASAP7_75t_R%SN VSS SN N_MM25_d N_MM16_s N_MM22_d N_MM15_d N_SN_11
+ N_SN_9 N_SN_10 N_SN_8 N_SN_12 N_SN_7 N_SN_1 N_SN_2 N_SN_15 N_SN_16
+ PM_FAx1_ASAP7_75t_R%SN
cc_109 N_SN_11 N_A_17 0.000179855f
cc_110 N_SN_11 N_MM21_g 0.000540252f
cc_111 N_SN_11 N_A_2 0.000349013f
cc_112 N_SN_9 N_A_2 0.000401242f
cc_113 N_SN_10 N_A_12 0.000460347f
cc_114 N_SN_9 N_A_17 0.000596238f
cc_115 N_SN_8 N_MM21_g 0.00106243f
cc_116 N_SN_12 N_A_17 0.00245059f
cc_117 N_SN_9 N_A_12 0.0030562f
cc_118 N_SN_11 N_A_15 0.00525746f
cc_119 N_SN_9 N_B_15 0.000161993f
cc_120 N_SN_9 N_MM20_g 0.000259332f
cc_121 N_SN_9 N_B_2 0.00129285f
cc_122 N_SN_12 N_B_15 0.000971935f
cc_123 N_SN_9 N_B_11 0.00642551f
cc_124 N_SN_7 N_CI_10 0.00103567f
cc_125 N_SN_8 N_MM22_g 0.0153611f
cc_126 N_SN_10 N_CI_10 0.000523924f
cc_127 N_SN_1 N_CI_2 0.000700593f
cc_128 N_SN_1 N_CI_10 0.00103048f
cc_129 N_SN_2 N_MM22_g 0.00117014f
cc_130 N_SN_1 N_MM22_g 0.00127616f
cc_131 N_SN_9 N_CI_16 0.00155025f
cc_132 N_SN_8 N_CI_2 0.0016436f
cc_133 N_SN_7 N_MM22_g 0.0533499f
cc_134 N_SN_7 N_CON_19 0.000208705f
cc_135 N_SN_7 N_CON_13 0.000237156f
cc_136 N_SN_7 N_CON_15 0.000309976f
cc_137 N_SN_7 N_CON_18 0.000377077f
cc_138 N_SN_8 N_MM15_g 0.0150352f
cc_139 N_SN_1 N_CON_15 0.000528299f
cc_140 N_SN_1 N_CON_1 0.000543474f
cc_141 N_SN_2 N_MM15_g 0.000874707f
cc_142 N_SN_10 N_CON_21 0.00108772f
cc_143 N_SN_1 N_MM15_g 0.00113595f
cc_144 N_SN_8 N_CON_1 0.00142628f
cc_145 N_SN_9 N_CON_13 0.00165557f
cc_146 N_SN_15 N_CON_19 0.0017783f
cc_147 N_SN_9 N_CON_21 0.00218773f
cc_148 N_SN_7 N_MM15_g 0.0520108f
x_PM_FAx1_ASAP7_75t_R%CON VSS CON N_MM15_g N_MM8_s N_MM7_s N_MM5_d N_MM1_d
+ N_CON_12 N_CON_10 N_CON_11 N_CON_13 N_CON_3 N_CON_4 N_CON_16 N_CON_17
+ N_CON_15 N_CON_21 N_CON_14 N_CON_18 N_CON_1 N_CON_20 N_CON_19
+ PM_FAx1_ASAP7_75t_R%CON
cc_149 N_CON_12 N_A_13 6.83506e-20
cc_150 N_CON_12 N_A_2 8.10998e-20
cc_151 N_CON_10 N_MM6_g 0.000676014f
cc_152 N_CON_11 N_MM6_g 8.25196e-20
cc_153 N_CON_13 N_A_11 9.1437e-20
cc_154 N_CON_12 N_A_14 0.000532921f
cc_155 N_CON_3 N_MM6_g 0.000139757f
cc_156 N_CON_4 N_MM6_g 0.000146408f
cc_157 N_CON_16 N_A_11 0.000151297f
cc_158 N_MM15_g N_MM21_g 0.000158421f
cc_159 N_CON_13 N_A_1 0.000218054f
cc_160 N_CON_12 N_A_1 0.00131914f
cc_161 N_CON_17 N_A_14 0.000511958f
cc_162 N_CON_15 N_A_17 0.000639792f
cc_163 N_CON_21 N_A_12 0.0013199f
cc_164 N_CON_14 N_A_17 0.00325218f
cc_165 N_CON_12 N_A_11 0.00424716f
cc_166 N_CON_10 N_B_11 5.72586e-20
cc_167 N_CON_10 N_B_2 7.51771e-20
cc_168 N_CON_10 N_B_14 8.92863e-20
cc_169 N_CON_13 N_B_2 0.000117638f
cc_170 N_CON_3 N_B_14 0.000194654f
cc_171 N_CON_4 N_B_14 0.000221114f
cc_172 N_CON_15 N_B_15 0.000374052f
cc_173 N_CON_13 N_B_11 0.000461988f
cc_174 N_CON_11 N_MM5_g 0.015914f
cc_175 N_CON_14 N_B_13 0.000647835f
cc_176 N_CON_3 N_B_1 0.000966511f
cc_177 N_CON_3 N_MM5_g 0.00110359f
cc_178 N_CON_4 N_MM5_g 0.00124361f
cc_179 N_CON_10 N_B_1 0.00184774f
cc_180 N_CON_13 N_B_14 0.00258211f
cc_181 N_CON_14 N_B_14 0.00263892f
cc_182 N_CON_12 N_B_13 0.00296202f
cc_183 N_CON_21 N_B_15 0.00384844f
cc_184 N_CON_10 N_MM5_g 0.0549871f
cc_185 N_CON_14 N_CI_12 0.000291289f
cc_186 N_CON_18 N_CI_10 0.00031528f
cc_187 N_CON_21 N_CI_14 0.000332713f
cc_188 N_CON_1 N_CI_3 0.000880776f
cc_189 N_CON_11 N_MM1_g 0.0155756f
cc_190 N_CON_20 N_CI_14 0.000467949f
cc_191 N_CON_21 N_CI_10 0.000527952f
cc_192 N_CON_19 N_CI_16 0.00053978f
cc_193 N_CON_21 N_CI_12 0.000604012f
cc_194 N_CON_3 N_CI_1 0.000646637f
cc_195 N_CON_4 N_MM1_g 0.000875874f
cc_196 N_CON_3 N_MM1_g 0.000887383f
cc_197 N_CON_1 N_CI_2 0.00242106f
cc_198 N_CON_13 N_CI_13 0.00115255f
cc_199 N_CON_13 N_CI_12 0.00140097f
cc_200 N_CON_11 N_CI_1 0.00151294f
cc_201 N_MM15_g N_MM14_g 0.0016772f
cc_202 N_CON_19 N_CI_14 0.00181678f
cc_203 N_CON_15 N_CI_10 0.00261566f
cc_204 N_CON_13 N_CI_11 0.00290133f
cc_205 N_MM15_g N_MM22_g 0.00491952f
cc_206 N_CON_21 N_CI_16 0.0250573f
cc_207 N_CON_10 N_MM1_g 0.0539637f
x_PM_FAx1_ASAP7_75t_R%CI VSS CI N_MM1_g N_MM22_g N_MM14_g N_CI_10 N_CI_14
+ N_CI_15 N_CI_3 N_CI_2 N_CI_16 N_CI_11 N_CI_13 N_CI_1 N_CI_12
+ PM_FAx1_ASAP7_75t_R%CI
cc_208 N_MM22_g N_A_17 0.000100177f
cc_209 N_MM22_g N_A_12 0.000140093f
cc_210 N_CI_10 N_A_15 0.000165112f
cc_211 N_CI_14 N_A_16 0.000220821f
cc_212 N_CI_14 N_A_13 0.00090478f
cc_213 N_CI_15 N_A_3 0.000392348f
cc_214 N_CI_3 N_A_3 0.0012283f
cc_215 N_CI_2 N_A_2 0.00271968f
cc_216 N_CI_16 N_A_17 0.00116994f
cc_217 N_CI_16 N_A_12 0.00126656f
cc_218 N_CI_15 N_A_13 0.00171087f
cc_219 N_CI_10 N_A_12 0.00231019f
cc_220 N_MM14_g N_MM17_g 0.00331056f
cc_221 N_MM22_g N_MM21_g 0.0070825f
cc_222 N_CI_16 N_MM20_g 0.000185149f
cc_223 N_CI_16 N_B_13 0.000110917f
cc_224 N_CI_15 N_B_15 0.000131806f
cc_225 N_CI_14 N_B_15 0.000830667f
cc_226 N_CI_10 N_B_15 0.000666522f
cc_227 N_CI_11 N_B_1 0.000396943f
cc_228 N_CI_13 N_B_2 0.000420894f
cc_229 N_CI_16 N_B_11 0.000457745f
cc_230 N_CI_1 N_B_2 0.000459953f
cc_231 N_CI_12 N_B_15 0.000514304f
cc_232 N_CI_1 N_B_1 0.00191722f
cc_233 N_CI_11 N_B_14 0.00105563f
cc_234 N_CI_12 N_B_14 0.00135779f
cc_235 N_MM1_g N_MM2_g 0.00166076f
cc_236 N_CI_13 N_B_11 0.00167833f
cc_237 N_MM1_g N_MM5_g 0.00495521f
cc_238 N_CI_16 N_B_15 0.0278348f
x_PM_FAx1_ASAP7_75t_R%B VSS B N_MM5_g N_MM2_g N_MM20_g N_MM18_g N_B_14 N_B_13
+ N_B_11 N_B_15 N_B_1 N_B_12 N_B_2 N_B_3 PM_FAx1_ASAP7_75t_R%B
cc_239 N_B_14 N_A_17 0.000112679f
cc_240 N_B_13 N_A_17 0.000631166f
cc_241 N_B_11 N_A_17 0.000629899f
cc_242 N_B_15 N_A_15 0.000458185f
cc_243 N_B_1 N_A_1 0.00182834f
cc_244 N_B_12 N_A_16 0.000241948f
cc_245 N_B_2 N_A_2 0.00208528f
cc_246 N_B_12 N_A_13 0.00286102f
cc_247 N_B_15 N_A_16 0.000384534f
cc_248 N_B_15 N_A_12 0.000691949f
cc_249 N_B_3 N_A_3 0.00153676f
cc_250 N_MM18_g N_MM17_g 0.00331642f
cc_251 N_MM20_g N_MM21_g 0.00694832f
cc_252 N_MM5_g N_MM6_g 0.00698163f
cc_253 N_B_15 N_A_17 0.0385576f
x_PM_FAx1_ASAP7_75t_R%A VSS A N_MM9_g N_MM6_g N_MM21_g N_MM17_g N_A_17 N_A_15
+ N_A_1 N_A_16 N_A_2 N_A_13 N_A_12 N_A_3 N_A_11 N_A_14 PM_FAx1_ASAP7_75t_R%A
*END of FAx1_ASAP7_75t_R.pxi
.ENDS
** Design:	HAxp5_ASAP7_75t_R
* Created:	"Fri Aug 17 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "HAxp5_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "HAxp5_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_HAxp5_ASAP7_75t_R%noxref_15 VSS 1
c1 1 VSS 0.00541283f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_12 VSS 1
c1 1 VSS 0.00460471f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_16 VSS 1
c1 1 VSS 0.00485715f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_17 VSS 1
c1 1 VSS 0.0047792f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_13 VSS 1
c1 1 VSS 0.0315616f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_14 VSS 1
c1 1 VSS 0.00624476f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%SN VSS 22 18 31 33 1 11 12 3 2 13 10 14 15
c1 1 VSS 0.00661791f
c2 2 VSS 0.00595617f
c3 3 VSS 0.0079179f
c4 10 VSS 0.00268371f
c5 11 VSS 0.00343478f
c6 12 VSS 0.00355787f
c7 13 VSS 0.0177619f
c8 14 VSS 0.00313331f
c9 15 VSS 0.00553671f
c10 16 VSS 0.00281395f
r1 33 32 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r2 11 32 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.2025 $X2=0.2845 $Y2=0.2025
r3 12 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.2025 $X2=0.4300 $Y2=0.2025
r4 31 12 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.2025 $X2=0.4175 $Y2=0.2025
r5 1 27 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.2160
+ $X2=0.2700 $Y2=0.2340
r6 3 13 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.2025
+ $X2=0.4320 $Y2=0.2340
r7 27 28 17.839 $w=1.3e-08 $l=7.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r8 25 28 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4185
+ $Y=0.2340 $X2=0.3465 $Y2=0.2340
r9 13 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4455 $Y2=0.2340
r10 13 25 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.2340 $X2=0.4185 $Y2=0.2340
r11 16 23 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.2340 $X2=0.4590 $Y2=0.2160
r12 16 24 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4590 $Y=0.2340 $X2=0.4455 $Y2=0.2340
r13 22 23 12.1259 $w=1.3e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1640 $X2=0.4590 $Y2=0.2160
r14 22 21 16.7897 $w=1.3e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.1640 $X2=0.4590 $Y2=0.0920
r15 14 20 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0360
r16 14 21 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4590
+ $Y=0.0540 $X2=0.4590 $Y2=0.0920
r17 19 20 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4455 $Y=0.0360 $X2=0.4590 $Y2=0.0360
r18 15 19 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.4320
+ $Y=0.0360 $X2=0.4455 $Y2=0.0360
r19 2 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.4320 $Y=0.0675
+ $X2=0.4320 $Y2=0.0360
r20 10 2 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4175 $Y=0.0675 $X2=0.4300 $Y2=0.0675
r21 18 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.4150 $Y=0.0675 $X2=0.4175 $Y2=0.0675
r22 1 11 1e-05
.ends

.subckt PM_HAxp5_ASAP7_75t_R%NET43 VSS 2 3 1
c1 1 VSS 0.000937793f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.1080 $Y2=0.0675
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.0675 $X2=0.1080 $Y2=0.0675
.ends

.subckt PM_HAxp5_ASAP7_75t_R%NET041 VSS 2 3 1
c1 1 VSS 0.00100786f
r1 2 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3070 $Y=0.2025 $X2=0.3240 $Y2=0.2025
r2 3 1 0.209877 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3410 $Y=0.2025 $X2=0.3240 $Y2=0.2025
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_10 VSS 1
c1 1 VSS 0.0419889f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%noxref_11 VSS 1
c1 1 VSS 0.0321379f
.ends

.subckt PM_HAxp5_ASAP7_75t_R%B VSS 21 3 4 1 6 7 5
c1 1 VSS 0.00868681f
c2 3 VSS 0.0355514f
c3 4 VSS 0.0461831f
c4 5 VSS 0.00371675f
c5 6 VSS 0.00347024f
c6 7 VSS 0.00368977f
r1 7 24 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1980 $X2=0.1350 $Y2=0.1665
r2 6 23 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0720 $X2=0.1350 $Y2=0.1035
r3 4 19 5.04173 $w=1.215e-07 $l=0 $layer=LIG $thickness=5.2e-08 $X=0.2970
+ $Y=0.1350 $X2=0.2970 $Y2=0.1350
r4 22 24 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1435 $X2=0.1350 $Y2=0.1665
r5 21 22 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1435
r6 21 5 1.98211 $w=1.3e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1265
r7 5 23 5.36336 $w=1.3e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1265 $X2=0.1350 $Y2=0.1035
r8 17 19 10.5547 $w=1.466e-08 $l=1.25e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2845 $Y=0.1350 $X2=0.2970 $Y2=0.1350
r9 16 17 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08 $X=0.2700
+ $Y=0.1350 $X2=0.2845 $Y2=0.1350
r10 15 16 96.7394 $w=9.3e-09 $l=4.15e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.2285 $Y=0.1350 $X2=0.2700 $Y2=0.1350
r11 14 15 97.9049 $w=9.3e-09 $l=4.2e-08 $layer=LIG $thickness=4.8e-08 $X=0.1865
+ $Y=0.1350 $X2=0.2285 $Y2=0.1350
r12 13 14 57.1112 $w=9.3e-09 $l=2.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1620 $Y=0.1350 $X2=0.1865 $Y2=0.1350
r13 12 13 33.8005 $w=9.3e-09 $l=1.45e-08 $layer=LIG $thickness=4.8e-08
+ $X=0.1475 $Y=0.1350 $X2=0.1620 $Y2=0.1350
r14 10 12 6.06403 $w=1.04167e-08 $l=3e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.1445 $Y=0.1350 $X2=0.1475 $Y2=0.1350
r15 9 10 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1445 $Y2=0.1350
r16 21 9 28.9687 $w=1.6e-08 $l=1.8e-08 $layer=V0LIG $X=0.1350 $Y=0.1350
+ $X2=0.1350 $Y2=0.1350
r17 1 9 4.49071 $w=1.6e-08 $l=9.5e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r18 1 11 1.40189 $w=1.265e-08 $l=1e-09 $layer=LIG $thickness=4.8e-08 $X=0.1255
+ $Y=0.1350 $X2=0.1245 $Y2=0.1350
r19 3 9 4.56902 $w=1.27053e-07 $l=0 $layer=LIG $thickness=5.22105e-08 $X=0.1350
+ $Y=0.1350 $X2=0.1350 $Y2=0.1350
r20 3 11 1.4802 $w=2.16633e-07 $l=1.05e-08 $layer=LIG $thickness=5.5619e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1245 $Y2=0.1350
r21 3 12 6.14234 $w=1.8346e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.1350 $Y=0.1350 $X2=0.1475 $Y2=0.1350
.ends

.subckt PM_HAxp5_ASAP7_75t_R%NET015 VSS 11 18 19 8 1 2 9 7
c1 1 VSS 0.00700334f
c2 2 VSS 0.00708434f
c3 7 VSS 0.00370621f
c4 8 VSS 0.00338558f
c5 9 VSS 0.0113856f
r1 19 17 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3950 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r2 2 17 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3780 $Y=0.0675 $X2=0.3925 $Y2=0.0675
r3 8 2 0.179012 $w=8.1e-08 $l=1.45e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3635 $Y=0.0675 $X2=0.3780 $Y2=0.0675
r4 18 8 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.3610 $Y=0.0675 $X2=0.3635 $Y2=0.0675
r5 2 15 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.3780 $Y=0.0675
+ $X2=0.3780 $Y2=0.0360
r6 14 15 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.3645
+ $Y=0.0360 $X2=0.3780 $Y2=0.0360
r7 13 14 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.3195
+ $Y=0.0360 $X2=0.3645 $Y2=0.0360
r8 12 13 11.5429 $w=1.3e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.2700
+ $Y=0.0360 $X2=0.3195 $Y2=0.0360
r9 9 12 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.2585
+ $Y=0.0360 $X2=0.2700 $Y2=0.0360
r10 1 12 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.2700 $Y=0.0675
+ $X2=0.2700 $Y2=0.0360
r11 11 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.2870 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r12 7 10 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.2720 $Y=0.0675 $X2=0.2845 $Y2=0.0675
r13 1 7 1e-05
.ends

.subckt PM_HAxp5_ASAP7_75t_R%A VSS 25 5 6 1 12 10 2 17 9 8 13 16 18
c1 1 VSS 0.00556504f
c2 2 VSS 0.00412908f
c3 5 VSS 0.0715445f
c4 6 VSS 0.0825557f
c5 7 VSS 0.00738397f
c6 8 VSS 0.0110454f
c7 9 VSS 0.018686f
c8 10 VSS 0.00205018f
c9 11 VSS 0.000355261f
c10 12 VSS 0.00415365f
c11 13 VSS 0.00347301f
c12 14 VSS 0.00472799f
c13 15 VSS 0.00187024f
c14 16 VSS 0.00293456f
c15 17 VSS 0.000415355f
c16 18 VSS 0.000834113f
r1 2 41 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.3510 $Y=0.1350
+ $X2=0.3510 $Y2=0.1350
r2 6 2 5.04045 $w=1.32911e-07 $l=0 $layer=LIG $thickness=5.24444e-08 $X=0.3510
+ $Y=0.1350 $X2=0.3510 $Y2=0.1350
r3 40 41 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1235 $X2=0.3510 $Y2=0.1350
r4 13 18 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.1010 $X2=0.3510 $Y2=0.0720
r5 13 40 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1010 $X2=0.3510 $Y2=0.1235
r6 18 39 10.4768 $w=1.38654e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3510 $Y=0.0720 $X2=0.2990 $Y2=0.0720
r7 12 17 4.22671 $w=1.43953e-08 $l=2.4683e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2405 $Y=0.0720 $X2=0.2160 $Y2=0.0690
r8 12 39 13.6416 $w=1.3e-08 $l=5.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.2405
+ $Y=0.0720 $X2=0.2990 $Y2=0.0720
r9 11 16 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0360
r10 11 17 2.71097 $w=1.5e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0540 $X2=0.2160 $Y2=0.0690
r11 16 37 3.59766 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.2160
+ $Y=0.0360 $X2=0.1935 $Y2=0.0360
r12 36 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0360 $X2=0.1935 $Y2=0.0360
r13 35 36 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.0360 $X2=0.1710 $Y2=0.0360
r14 34 35 6.52931 $w=1.3e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1250
+ $Y=0.0360 $X2=0.1530 $Y2=0.0360
r15 33 34 5.82974 $w=1.3e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1000
+ $Y=0.0360 $X2=0.1250 $Y2=0.0360
r16 32 33 3.26466 $w=1.3e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.0860
+ $Y=0.0360 $X2=0.1000 $Y2=0.0360
r17 9 14 5.34658 $w=1.45e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.0360 $X2=0.0270 $Y2=0.0360
r18 9 32 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0570
+ $Y=0.0360 $X2=0.0860 $Y2=0.0360
r19 14 28 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0360 $X2=0.0270 $Y2=0.0540
r20 8 15 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1665 $X2=0.0270 $Y2=0.1350
r21 27 28 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0720 $X2=0.0270 $Y2=0.0540
r22 7 15 6.16517 $w=1.44286e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1035 $X2=0.0270 $Y2=0.1350
r23 7 27 7.34548 $w=1.3e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1035 $X2=0.0270 $Y2=0.0720
r24 25 10 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.0640
+ $Y=0.1350 $X2=0.0455 $Y2=0.1350
r25 10 15 3.1337 $w=1.54324e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0455 $Y=0.1350 $X2=0.0270 $Y2=0.1350
r26 25 23 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0640 $Y=0.1350
+ $X2=0.0605 $Y2=0.1350
r27 21 23 4.72579 $w=1.53e-08 $l=8e-09 $layer=LIG $thickness=4.8e-08 $X=0.0685
+ $Y=0.1350 $X2=0.0605 $Y2=0.1350
r28 1 20 2.6116 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=4.8e-08 $X=0.0720
+ $Y=0.1350 $X2=0.0820 $Y2=0.1350
r29 1 21 1.73797 $w=1.72143e-08 $l=3.5e-09 $layer=LIG $thickness=4.8e-08
+ $X=0.0720 $Y=0.1350 $X2=0.0685 $Y2=0.1350
r30 5 20 2.66511 $w=1.29895e-07 $l=1e-09 $layer=LIG $thickness=5.22105e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0820 $Y2=0.1350
r31 5 21 1.79147 $w=1.8466e-07 $l=1.25e-08 $layer=LIG $thickness=5.44e-08
+ $X=0.0810 $Y=0.1350 $X2=0.0685 $Y2=0.1350
.ends

.subckt PM_HAxp5_ASAP7_75t_R%CON VSS 27 9 35 43 44 13 11 4 3 12 1 15 16 10 14
+ 17 19
c1 1 VSS 0.00167818f
c2 3 VSS 0.0088938f
c3 4 VSS 0.00619887f
c4 9 VSS 0.0421499f
c5 10 VSS 0.00468381f
c6 11 VSS 0.00581189f
c7 12 VSS 0.00723799f
c8 13 VSS 0.00191503f
c9 14 VSS 0.000786088f
c10 15 VSS 0.00681414f
c11 16 VSS 0.00157385f
c12 17 VSS 0.000512191f
c13 18 VSS 0.00274833f
c14 19 VSS 0.000425887f
r1 44 42 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.1250 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r2 3 42 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1080 $Y=0.2160 $X2=0.1225 $Y2=0.2160
r3 11 3 0.268519 $w=5.4e-08 $l=1.45e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2160 $X2=0.1080 $Y2=0.2160
r4 43 11 0.0462963 $w=5.4e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2160 $X2=0.0935 $Y2=0.2160
r5 3 36 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2160
+ $X2=0.1120 $Y2=0.2340
r6 36 37 4.31401 $w=1.3e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.1120
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r7 12 18 2.5483 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1710 $Y2=0.2340
r8 12 37 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1530
+ $Y=0.2340 $X2=0.1305 $Y2=0.2340
r9 10 4 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1475 $Y=0.0675 $X2=0.1600 $Y2=0.0675
r10 35 10 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.1450 $Y=0.0675 $X2=0.1475 $Y2=0.0675
r11 4 31 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1745 $Y=0.0675
+ $X2=0.1710 $Y2=0.0900
r12 14 17 3.01711 $w=1.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.2160 $X2=0.1710 $Y2=0.1980
r13 14 18 2.5483 $w=1.79e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.2160 $X2=0.1710 $Y2=0.2340
r14 31 32 8.04505 $w=1.3e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.0900 $X2=0.1710 $Y2=0.1245
r15 13 17 5.4656 $w=1.45789e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1710 $Y=0.1695 $X2=0.1710 $Y2=0.1980
r16 13 32 10.4935 $w=1.3e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1695 $X2=0.1710 $Y2=0.1245
r17 17 30 4.06646 $w=1.5e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1710
+ $Y=0.1980 $X2=0.1935 $Y2=0.1980
r18 29 30 8.86121 $w=1.3e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2315
+ $Y=0.1980 $X2=0.1935 $Y2=0.1980
r19 27 28 9.96886 $w=1.3e-08 $l=4.27e-08 $layer=M1 $thickness=3.6e-08 $X=0.2570
+ $Y=0.1980 $X2=0.2997 $Y2=0.1980
r20 27 26 0.174892 $w=1.3e-08 $l=8e-10 $layer=M1 $thickness=3.6e-08 $X=0.2570
+ $Y=0.1980 $X2=0.2562 $Y2=0.1980
r21 26 29 5.77145 $w=1.3e-08 $l=2.47e-08 $layer=M1 $thickness=3.6e-08 $X=0.2562
+ $Y=0.1980 $X2=0.2315 $Y2=0.1980
r22 25 28 11.951 $w=1.3e-08 $l=5.13e-08 $layer=M1 $thickness=3.6e-08 $X=0.3510
+ $Y=0.1980 $X2=0.2997 $Y2=0.1980
r23 24 25 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.3735
+ $Y=0.1980 $X2=0.3510 $Y2=0.1980
r24 15 19 1.49895 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.3915 $Y=0.1980 $X2=0.4050 $Y2=0.1980
r25 15 24 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.3915
+ $Y=0.1980 $X2=0.3735 $Y2=0.1980
r26 19 23 4.9968 $w=1.60947e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4050 $Y=0.1980 $X2=0.4050 $Y2=0.1695
r27 22 23 5.24677 $w=1.3e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1470 $X2=0.4050 $Y2=0.1695
r28 21 22 2.79828 $w=1.3e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1470
r29 16 21 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.4050
+ $Y=0.1235 $X2=0.4050 $Y2=0.1350
r30 9 1 6.81262 $w=1.1611e-07 $l=0 $layer=LIG $thickness=5.18095e-08 $X=0.4050
+ $Y=0.1350 $X2=0.4050 $Y2=0.1350
r31 1 21 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.4050 $Y=0.1350
+ $X2=0.4050 $Y2=0.1350
.ends


*
.SUBCKT HAxp5_ASAP7_75t_R VSS VDD A B CON SN
*
* VSS VSS
* VDD VDD
* A A
* B B
* CON CON
* SN SN
*
*

MM3 N_MM3_d N_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM2 N_MM2_d N_MM2_g N_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM5 N_MM5_d N_MM5_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM4 N_MM4_d N_MM4_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM6 N_MM6_d N_MM6_g N_MM6_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM0 N_MM0_d N_MM3_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM1 N_MM1_d N_MM2_g VDD VDD pmos_rvt L=2e-08 W=5.4e-08 nfin=2
MM10 N_MM10_d N_MM5_g N_MM10_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM11 N_MM11_d N_MM4_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM9 N_MM9_d N_MM6_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "HAxp5_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "HAxp5_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_HAxp5_ASAP7_75t_R%noxref_15 VSS N_noxref_15_1
+ PM_HAxp5_ASAP7_75t_R%noxref_15
cc_1 N_noxref_15_1 N_B_1 0.00113715f
cc_2 N_noxref_15_1 N_MM5_g 0.0023561f
cc_3 N_noxref_15_1 N_SN_11 0.0365475f
cc_4 N_noxref_15_1 N_noxref_13_1 0.00749033f
cc_5 N_noxref_15_1 N_noxref_14_1 0.000895268f
x_PM_HAxp5_ASAP7_75t_R%noxref_12 VSS N_noxref_12_1
+ PM_HAxp5_ASAP7_75t_R%noxref_12
cc_6 N_noxref_12_1 N_B_1 0.000991179f
cc_7 N_noxref_12_1 N_MM2_g 0.00228133f
cc_8 N_noxref_12_1 N_CON_4 0.00158701f
cc_9 N_noxref_12_1 N_CON_10 0.0368277f
x_PM_HAxp5_ASAP7_75t_R%noxref_16 VSS N_noxref_16_1
+ PM_HAxp5_ASAP7_75t_R%noxref_16
cc_10 N_noxref_16_1 N_MM6_g 0.00145624f
cc_11 N_noxref_16_1 N_SN_10 0.0383353f
x_PM_HAxp5_ASAP7_75t_R%noxref_17 VSS N_noxref_17_1
+ PM_HAxp5_ASAP7_75t_R%noxref_17
cc_12 N_noxref_17_1 N_MM6_g 0.00145722f
cc_13 N_noxref_17_1 N_SN_12 0.0384726f
cc_14 N_noxref_17_1 N_noxref_16_1 0.00177384f
x_PM_HAxp5_ASAP7_75t_R%noxref_13 VSS N_noxref_13_1
+ PM_HAxp5_ASAP7_75t_R%noxref_13
cc_15 N_noxref_13_1 N_B_1 0.00138916f
cc_16 N_noxref_13_1 N_MM2_g 0.00431442f
cc_17 N_noxref_13_1 N_CON_11 0.000512876f
cc_18 N_noxref_13_1 N_noxref_12_1 0.000965398f
x_PM_HAxp5_ASAP7_75t_R%noxref_14 VSS N_noxref_14_1
+ PM_HAxp5_ASAP7_75t_R%noxref_14
cc_19 N_noxref_14_1 N_B_1 0.00108047f
cc_20 N_noxref_14_1 N_MM5_g 0.00230394f
cc_21 N_noxref_14_1 N_CON_4 0.00100694f
cc_22 N_noxref_14_1 N_NET015_7 0.0351074f
cc_23 N_noxref_14_1 N_noxref_12_1 0.00731502f
x_PM_HAxp5_ASAP7_75t_R%SN VSS SN N_MM6_d N_MM9_d N_MM10_d N_SN_1 N_SN_11
+ N_SN_12 N_SN_3 N_SN_2 N_SN_13 N_SN_10 N_SN_14 N_SN_15 PM_HAxp5_ASAP7_75t_R%SN
cc_24 N_SN_1 N_MM5_g 0.0018131f
cc_25 N_SN_11 N_B_1 0.0023775f
cc_26 N_SN_11 N_MM5_g 0.0359805f
cc_27 N_SN_12 N_MM6_g 0.0158483f
cc_28 N_SN_3 N_CON_1 0.00085171f
cc_29 N_SN_2 N_MM6_g 0.00107049f
cc_30 N_SN_1 N_CON_15 0.00121726f
cc_31 N_SN_3 N_MM6_g 0.00140523f
cc_32 N_SN_13 N_CON_19 0.00145328f
cc_33 N_SN_10 N_CON_1 0.00157844f
cc_34 N_SN_14 N_CON_16 0.00447808f
cc_35 N_SN_13 N_CON_15 0.0136874f
cc_36 N_SN_10 N_MM6_g 0.0547139f
cc_37 N_SN_15 N_NET015_9 0.00074869f
cc_38 N_SN_2 N_NET015_2 0.00516316f
x_PM_HAxp5_ASAP7_75t_R%NET43 VSS N_MM3_d N_MM2_s N_NET43_1
+ PM_HAxp5_ASAP7_75t_R%NET43
cc_39 N_NET43_1 N_MM3_g 0.0174944f
cc_40 N_NET43_1 N_MM2_g 0.0174018f
x_PM_HAxp5_ASAP7_75t_R%NET041 VSS N_MM10_s N_MM11_d N_NET041_1
+ PM_HAxp5_ASAP7_75t_R%NET041
cc_41 N_NET041_1 N_MM4_g 0.0172237f
cc_42 N_NET041_1 N_MM5_g 0.0174148f
x_PM_HAxp5_ASAP7_75t_R%noxref_10 VSS N_noxref_10_1
+ PM_HAxp5_ASAP7_75t_R%noxref_10
cc_43 N_noxref_10_1 N_MM3_g 0.00263963f
x_PM_HAxp5_ASAP7_75t_R%noxref_11 VSS N_noxref_11_1
+ PM_HAxp5_ASAP7_75t_R%noxref_11
cc_44 N_noxref_11_1 N_MM3_g 0.00466932f
cc_45 N_noxref_11_1 N_noxref_10_1 0.00185044f
x_PM_HAxp5_ASAP7_75t_R%B VSS B N_MM2_g N_MM5_g N_B_1 N_B_6 N_B_7 N_B_5
+ PM_HAxp5_ASAP7_75t_R%B
cc_46 N_B_1 N_MM3_g 0.000368993f
cc_47 N_B_6 N_MM3_g 0.000272835f
cc_48 N_B_7 N_MM3_g 0.000327878f
cc_49 N_B_1 N_A_1 0.00179117f
cc_50 N_B_1 N_A_12 0.000424587f
cc_51 N_B_7 N_A_10 0.000480064f
cc_52 N_B_1 N_A_2 0.000487389f
cc_53 N_B_1 N_A_17 0.00196061f
cc_54 N_B_5 N_A_10 0.00216126f
cc_55 N_B_6 N_A_9 0.00482503f
cc_56 N_MM5_g N_MM4_g 0.00490939f
cc_57 N_MM2_g N_MM3_g 0.00743415f
x_PM_HAxp5_ASAP7_75t_R%NET015 VSS N_MM5_d N_MM4_d N_MM6_s N_NET015_8 N_NET015_1
+ N_NET015_2 N_NET015_9 N_NET015_7 PM_HAxp5_ASAP7_75t_R%NET015
cc_58 N_NET015_8 N_A_16 0.000475473f
cc_59 N_NET015_1 N_A_12 0.00156071f
cc_60 N_NET015_2 N_A_13 0.000600565f
cc_61 N_NET015_8 N_A_2 0.000778719f
cc_62 N_NET015_2 N_MM4_g 0.00129272f
cc_63 N_NET015_9 N_A_18 0.001342f
cc_64 N_NET015_9 N_A_12 0.0084283f
cc_65 N_NET015_8 N_MM4_g 0.0341513f
cc_66 N_NET015_1 N_MM5_g 0.00154348f
cc_67 N_NET015_7 N_B_1 0.00212346f
cc_68 N_NET015_7 N_MM5_g 0.0339689f
cc_69 N_NET015_8 N_CON_4 0.000422117f
cc_70 N_NET015_7 N_CON_4 0.000578916f
cc_71 N_NET015_8 N_CON_1 0.000663398f
cc_72 N_NET015_2 N_MM6_g 0.00090459f
cc_73 N_NET015_8 N_MM6_g 0.0340905f
x_PM_HAxp5_ASAP7_75t_R%A VSS A N_MM3_g N_MM4_g N_A_1 N_A_12 N_A_10 N_A_2 N_A_17
+ N_A_9 N_A_8 N_A_13 N_A_16 N_A_18 PM_HAxp5_ASAP7_75t_R%A
x_PM_HAxp5_ASAP7_75t_R%CON VSS CON N_MM6_g N_MM2_d N_MM0_d N_MM1_d N_CON_13
+ N_CON_11 N_CON_4 N_CON_3 N_CON_12 N_CON_1 N_CON_15 N_CON_16 N_CON_10 N_CON_14
+ N_CON_17 N_CON_19 PM_HAxp5_ASAP7_75t_R%CON
cc_74 N_CON_13 N_MM3_g 0.000292027f
cc_75 N_CON_11 N_A_1 0.000369571f
cc_76 N_CON_4 N_A_17 0.000498853f
cc_77 N_CON_3 N_MM3_g 0.000610858f
cc_78 N_CON_12 N_A_8 0.000769181f
cc_79 N_CON_4 N_A_12 0.00079663f
cc_80 N_CON_1 N_A_2 0.00198511f
cc_81 N_CON_15 N_A_13 0.00162059f
cc_82 N_CON_4 N_A_9 0.00163508f
cc_83 N_CON_13 N_A_9 0.00167388f
cc_84 N_CON_13 N_A_17 0.00260546f
cc_85 N_CON_16 N_A_13 0.00293113f
cc_86 N_MM6_g N_MM4_g 0.00338312f
cc_87 N_CON_11 N_MM3_g 0.0263953f
cc_88 N_CON_10 N_B_7 0.000252713f
cc_89 N_CON_14 N_B_7 0.000402489f
cc_90 N_CON_13 N_B_1 0.000724088f
cc_91 N_CON_4 N_B_5 0.00075426f
cc_92 N_CON_3 N_MM2_g 0.000845936f
cc_93 N_CON_13 N_B_6 0.000856128f
cc_94 N_CON_15 N_B_1 0.000927972f
cc_95 N_CON_17 N_B_7 0.00261946f
cc_96 N_CON_4 N_MM2_g 0.00315994f
cc_97 N_CON_12 N_B_7 0.00328825f
cc_98 N_CON_11 N_MM2_g 0.0109967f
cc_99 N_CON_4 N_B_1 0.00488079f
cc_100 N_CON_13 N_B_5 0.00988383f
cc_101 N_CON_10 N_MM2_g 0.0500158f
*END of HAxp5_ASAP7_75t_R.pxi
.ENDS
** Design:	TIEHIx1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "TIEHIx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "TIEHIx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_TIEHIx1_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.0200419f
.ends

.subckt PM_TIEHIx1_ASAP7_75t_R%noxref_5 VSS 1
c1 1 VSS 0.00429921f
.ends

.subckt PM_TIEHIx1_ASAP7_75t_R%noxref_6 VSS 1
c1 1 VSS 0.0431249f
.ends

.subckt PM_TIEHIx1_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.00502181f
.ends

.subckt PM_TIEHIx1_ASAP7_75t_R%NET7 VSS 6 28 3 1 8 9 10 7
c1 1 VSS 0.00406377f
c2 3 VSS 0.00633118f
c3 6 VSS 0.0400772f
c4 7 VSS 0.00379302f
c5 8 VSS 0.00420362f
c6 9 VSS 0.0023873f
c7 10 VSS 0.00752476f
c8 11 VSS 0.00189164f
r1 28 27 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.0405 $X2=0.0685 $Y2=0.0405
r2 7 27 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.0405 $X2=0.0685 $Y2=0.0405
r3 3 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.0405
+ $X2=0.0540 $Y2=0.0360
r4 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.0360 $X2=0.0540 $Y2=0.0360
r5 10 22 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0270 $Y2=0.0575
r6 10 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.0360 $X2=0.0405 $Y2=0.0360
r7 21 22 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.0790 $X2=0.0270 $Y2=0.0575
r8 8 11 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1080 $X2=0.0270 $Y2=0.1370
r9 8 21 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1080 $X2=0.0270 $Y2=0.0790
r10 11 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1370 $X2=0.0515 $Y2=0.1370
r11 9 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1370 $X2=0.0810 $Y2=0.1370
r12 9 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1370 $X2=0.0515 $Y2=0.1370
r13 1 12 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1370 $X2=0.0810 $Y2=0.1370
r14 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1370
+ $X2=0.0810 $Y2=0.1370
r15 6 12 0.558039 $w=1.28e-07 $l=4.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.1845 $X2=0.0810 $Y2=0.1370
r16 3 7 1e-05
.ends

.subckt PM_TIEHIx1_ASAP7_75t_R%H VSS 23 6 30 1 3 8 9 7
c1 1 VSS 0.00448065f
c2 3 VSS 0.0088639f
c3 6 VSS 0.0180104f
c4 7 VSS 0.00443935f
c5 8 VSS 0.00193559f
c6 9 VSS 0.00436299f
c7 10 VSS 0.00666584f
c8 11 VSS 0.00159257f
r1 7 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.2025 $X2=0.1060 $Y2=0.2025
r2 30 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.2025 $X2=0.0935 $Y2=0.2025
r3 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.2025
+ $X2=0.1080 $Y2=0.2340
r4 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.2340 $X2=0.1215 $Y2=0.2340
r5 10 24 4.53284 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.2340 $X2=0.1350 $Y2=0.2095
r6 10 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.2340 $X2=0.1215 $Y2=0.2340
r7 23 24 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1935 $X2=0.1350 $Y2=0.2095
r8 23 22 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1935 $X2=0.1350 $Y2=0.1695
r9 21 22 7.57867 $w=1.3e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1370 $X2=0.1350 $Y2=0.1695
r10 9 11 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1080 $X2=0.1350 $Y2=0.0790
r11 9 21 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1080 $X2=0.1350 $Y2=0.1370
r12 11 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0790 $X2=0.1105 $Y2=0.0790
r13 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0925
+ $Y=0.0790 $X2=0.1105 $Y2=0.0790
r14 18 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.0790 $X2=0.0925 $Y2=0.0790
r15 17 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.0790 $X2=0.0810 $Y2=0.0790
r16 8 17 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.0790 $X2=0.0700 $Y2=0.0790
r17 1 12 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.0790 $X2=0.0810 $Y2=0.0790
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.0790
+ $X2=0.0810 $Y2=0.0790
r19 6 12 0.860591 $w=8.3e-08 $l=1.6e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.0630 $X2=0.0810 $Y2=0.0790
.ends


*
.SUBCKT TIEHIx1_ASAP7_75t_R VSS VDD H
*
* VSS VSS
* VDD VDD
* H H
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=2.7e-08 nfin=1
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3


*include "TIEHIx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "TIEHIx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_TIEHIx1_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_TIEHIx1_ASAP7_75t_R%noxref_7
cc_1 N_noxref_7_1 N_MM2_g 0.00145024f
cc_2 N_noxref_7_1 N_H_1 0.00345257f
cc_3 N_noxref_7_1 N_NET7_7 0.000929614f
x_PM_TIEHIx1_ASAP7_75t_R%noxref_5 VSS N_noxref_5_1
+ PM_TIEHIx1_ASAP7_75t_R%noxref_5
cc_4 N_noxref_5_1 N_H_1 0.00411826f
cc_5 N_noxref_5_1 N_NET7_7 0.0177076f
x_PM_TIEHIx1_ASAP7_75t_R%noxref_6 VSS N_noxref_6_1
+ PM_TIEHIx1_ASAP7_75t_R%noxref_6
cc_6 N_noxref_6_1 N_H_7 0.000901816f
cc_7 N_noxref_6_1 N_MM1_g 0.00430527f
cc_8 N_noxref_6_1 N_noxref_5_1 0.00602471f
x_PM_TIEHIx1_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_TIEHIx1_ASAP7_75t_R%noxref_8
cc_9 N_noxref_8_1 N_H_7 0.0399543f
cc_10 N_noxref_8_1 N_MM1_g 0.00353069f
cc_11 N_noxref_8_1 N_noxref_7_1 0.00602361f
x_PM_TIEHIx1_ASAP7_75t_R%NET7 VSS N_MM1_g N_MM2_d N_NET7_3 N_NET7_1 N_NET7_8
+ N_NET7_9 N_NET7_10 N_NET7_7 PM_TIEHIx1_ASAP7_75t_R%NET7
cc_12 N_NET7_3 N_H_1 0.00250407f
cc_13 N_NET7_1 N_H_3 0.000968018f
cc_14 N_NET7_8 N_H_8 0.00141865f
cc_15 N_MM1_g N_H_3 0.00153513f
cc_16 N_NET7_9 N_H_9 0.00178819f
cc_17 N_NET7_9 N_H_8 0.00198057f
cc_18 N_NET7_10 N_H_8 0.00296245f
cc_19 N_NET7_1 N_H_7 0.00322065f
cc_20 N_NET7_7 N_H_1 0.00338016f
cc_21 N_NET7_7 N_MM2_g 0.0177435f
cc_22 N_MM1_g N_H_7 0.0383611f
x_PM_TIEHIx1_ASAP7_75t_R%H VSS H N_MM2_g N_MM1_d N_H_1 N_H_3 N_H_8 N_H_9 N_H_7
+ PM_TIEHIx1_ASAP7_75t_R%H
*END of TIEHIx1_ASAP7_75t_R.pxi
.ENDS
** Design:	TIELOx1_ASAP7_75t_R
* Created:	"Sat Aug 18 2018"
* Vendor:	"Mentor Graphics Corporation"
* Program:	"xACT"
* Version:	"v2017.1_34.33"
* Corner Name: typical_27
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* Integrated TICER reduction is not enabled.
* SHORT DELAY THRESHOLD: 2e-15
* Fill Mode: NG
* PEX REDUCE CC ABSOLUTE : 1
* PEX REDUCE CC RELATIVE : 0.01
* Delta transform mode : 344834

*include "TIELOx1_ASAP7_75t_R.pex.netlist.pex"
*BEGIN of ".include "TIELOx1_ASAP7_75t_R.pex.netlist.pex"


.subckt PM_TIELOx1_ASAP7_75t_R%noxref_5 VSS 1
c1 1 VSS 0.0431249f
.ends

.subckt PM_TIELOx1_ASAP7_75t_R%noxref_6 VSS 1
c1 1 VSS 0.00429921f
.ends

.subckt PM_TIELOx1_ASAP7_75t_R%noxref_7 VSS 1
c1 1 VSS 0.00502264f
.ends

.subckt PM_TIELOx1_ASAP7_75t_R%NET9 VSS 6 28 3 1 8 9 11 7
c1 1 VSS 0.00406365f
c2 3 VSS 0.00633103f
c3 6 VSS 0.0400772f
c4 7 VSS 0.00379207f
c5 8 VSS 0.00420166f
c6 9 VSS 0.00238642f
c7 10 VSS 0.00189083f
c8 11 VSS 0.00752386f
r1 28 27 0.0925926 $w=2.7e-08 $l=2.5e-09 $layer=P_src_drn $thickness=1e-09
+ $X=0.0710 $Y=0.2295 $X2=0.0685 $Y2=0.2295
r2 7 27 0.462963 $w=2.7e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.0560 $Y=0.2295 $X2=0.0685 $Y2=0.2295
r3 3 24 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.0540 $Y=0.2295
+ $X2=0.0540 $Y2=0.2340
r4 23 24 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.0405
+ $Y=0.2340 $X2=0.0540 $Y2=0.2340
r5 11 22 3.83327 $w=1.5093e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0270 $Y2=0.2125
r6 11 23 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.2340 $X2=0.0405 $Y2=0.2340
r7 21 22 5.01358 $w=1.3e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1910 $X2=0.0270 $Y2=0.2125
r8 8 10 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1620 $X2=0.0270 $Y2=0.1330
r9 8 21 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.0270
+ $Y=0.1620 $X2=0.0270 $Y2=0.1910
r10 10 19 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.0270 $Y=0.1330 $X2=0.0515 $Y2=0.1330
r11 9 17 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1330 $X2=0.0810 $Y2=0.1330
r12 9 19 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0695
+ $Y=0.1330 $X2=0.0515 $Y2=0.1330
r13 1 12 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1330 $X2=0.0810 $Y2=0.1330
r14 1 17 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1330
+ $X2=0.0810 $Y2=0.1330
r15 6 12 0.558039 $w=1.28e-07 $l=4.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.0855 $X2=0.0810 $Y2=0.1330
r16 3 7 1e-05
.ends

.subckt PM_TIELOx1_ASAP7_75t_R%noxref_8 VSS 1
c1 1 VSS 0.0200419f
.ends

.subckt PM_TIELOx1_ASAP7_75t_R%L VSS 23 6 30 1 3 8 9 7
c1 1 VSS 0.00448098f
c2 3 VSS 0.00886514f
c3 6 VSS 0.0180104f
c4 7 VSS 0.00444459f
c5 8 VSS 0.00193772f
c6 9 VSS 0.00437302f
c7 10 VSS 0.0070593f
c8 11 VSS 0.00159473f
r1 7 3 0.154321 $w=8.1e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.0935 $Y=0.0675 $X2=0.1060 $Y2=0.0675
r2 30 7 0.0308642 $w=8.1e-08 $l=2.5e-09 $layer=N_src_drn $thickness=1e-09
+ $X=0.0910 $Y=0.0675 $X2=0.0935 $Y2=0.0675
r3 3 26 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LISD $X=0.1080 $Y=0.0675
+ $X2=0.1080 $Y2=0.0360
r4 26 27 3.14806 $w=1.3e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.1080
+ $Y=0.0360 $X2=0.1215 $Y2=0.0360
r5 10 22 4.53284 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0360 $X2=0.1350 $Y2=0.0605
r6 10 27 1.96775 $w=1.63333e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.0360 $X2=0.1215 $Y2=0.0360
r7 23 24 5.59655 $w=1.3e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0765 $X2=0.1350 $Y2=0.1005
r8 23 22 3.73104 $w=1.3e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.0765 $X2=0.1350 $Y2=0.0605
r9 21 24 7.57867 $w=1.3e-08 $l=3.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1330 $X2=0.1350 $Y2=0.1005
r10 9 11 5.11339 $w=1.60414e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1620 $X2=0.1350 $Y2=0.1910
r11 9 21 6.7625 $w=1.3e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.1350
+ $Y=0.1620 $X2=0.1350 $Y2=0.1330
r12 11 20 4.06404 $w=1.48367e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.1350 $Y=0.1910 $X2=0.1105 $Y2=0.1910
r13 19 20 4.19742 $w=1.3e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.0925
+ $Y=0.1910 $X2=0.1105 $Y2=0.1910
r14 18 19 2.68168 $w=1.3e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.0810
+ $Y=0.1910 $X2=0.0925 $Y2=0.1910
r15 17 18 2.56509 $w=1.3e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.0700
+ $Y=0.1910 $X2=0.0810 $Y2=0.1910
r16 8 17 0.582974 $w=1.3e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0675
+ $Y=0.1910 $X2=0.0700 $Y2=0.1910
r17 1 12 2.6116 $w=2.2e-08 $l=0 $layer=LIG $thickness=4.8e-08 $X=0.0810
+ $Y=0.1910 $X2=0.0810 $Y2=0.1910
r18 1 18 19.3796 $w=1.8e-08 $l=1.8e-08 $layer=V0LIG $X=0.0810 $Y=0.1910
+ $X2=0.0810 $Y2=0.1910
r19 6 12 0.860591 $w=8.3e-08 $l=1.6e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.0810 $Y=0.2070 $X2=0.0810 $Y2=0.1910
.ends


*
.SUBCKT TIELOx1_ASAP7_75t_R VSS VDD L
*
* VSS VSS
* VDD VDD
* L L
*
*

MM2 N_MM2_d N_MM2_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
MM1 N_MM1_d N_MM1_g VDD VDD pmos_rvt L=2e-08 W=2.7e-08 nfin=1


*include "TIELOx1_ASAP7_75t_R.pex.netlist.pxi"
*BEGIN of ".include "TIELOx1_ASAP7_75t_R.pex.netlist.pxi"

*ENDS
*
x_PM_TIELOx1_ASAP7_75t_R%noxref_5 VSS N_noxref_5_1
+ PM_TIELOx1_ASAP7_75t_R%noxref_5
cc_1 N_noxref_5_1 N_MM2_g 0.00430527f
cc_2 N_noxref_5_1 N_L_7 0.000901816f
x_PM_TIELOx1_ASAP7_75t_R%noxref_6 VSS N_noxref_6_1
+ PM_TIELOx1_ASAP7_75t_R%noxref_6
cc_3 N_noxref_6_1 N_NET9_7 0.0177076f
cc_4 N_noxref_6_1 N_L_1 0.00411826f
cc_5 N_noxref_6_1 N_noxref_5_1 0.00602471f
x_PM_TIELOx1_ASAP7_75t_R%noxref_7 VSS N_noxref_7_1
+ PM_TIELOx1_ASAP7_75t_R%noxref_7
cc_6 N_noxref_7_1 N_MM2_g 0.00353069f
cc_7 N_noxref_7_1 N_L_7 0.0399535f
x_PM_TIELOx1_ASAP7_75t_R%NET9 VSS N_MM2_g N_MM1_d N_NET9_3 N_NET9_1 N_NET9_8
+ N_NET9_9 N_NET9_11 N_NET9_7 PM_TIELOx1_ASAP7_75t_R%NET9
x_PM_TIELOx1_ASAP7_75t_R%noxref_8 VSS N_noxref_8_1
+ PM_TIELOx1_ASAP7_75t_R%noxref_8
cc_8 N_noxref_8_1 N_NET9_7 0.000929614f
cc_9 N_noxref_8_1 N_MM1_g 0.00145024f
cc_10 N_noxref_8_1 N_L_1 0.00345272f
cc_11 N_noxref_8_1 N_noxref_7_1 0.00602361f
x_PM_TIELOx1_ASAP7_75t_R%L VSS L N_MM1_g N_MM2_d N_L_1 N_L_3 N_L_8 N_L_9 N_L_7
+ PM_TIELOx1_ASAP7_75t_R%L
cc_12 N_L_1 N_NET9_3 0.00250407f
cc_13 N_L_3 N_NET9_1 0.000968018f
cc_14 N_L_8 N_NET9_8 0.00141865f
cc_15 N_L_3 N_MM2_g 0.00153513f
cc_16 N_L_9 N_NET9_9 0.00178819f
cc_17 N_L_8 N_NET9_9 0.00198057f
cc_18 N_L_8 N_NET9_11 0.00296245f
cc_19 N_L_7 N_NET9_1 0.00322065f
cc_20 N_L_1 N_NET9_7 0.00338016f
cc_21 N_MM1_g N_NET9_7 0.0177435f
cc_22 N_L_7 N_MM2_g 0.0383669f
*END of TIELOx1_ASAP7_75t_R.pxi
.ENDS
*